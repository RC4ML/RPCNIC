module MMCME4_ADV_Wrapper(
  input   io_CLKIN1,
  output  io_LOCKED,
  output  io_CLKOUT0,
  output  io_CLKOUT1,
  output  io_CLKOUT2,
  output  io_CLKOUT3,
  output  io_CLKOUT4,
  output  io_CLKOUT5
);
  wire  mmcm4_adv_CLKIN1; // @[Buf.scala 109:25]
  wire  mmcm4_adv_CLKIN2; // @[Buf.scala 109:25]
  wire  mmcm4_adv_RST; // @[Buf.scala 109:25]
  wire  mmcm4_adv_PWRDWN; // @[Buf.scala 109:25]
  wire  mmcm4_adv_CDDCREQ; // @[Buf.scala 109:25]
  wire  mmcm4_adv_CLKINSEL; // @[Buf.scala 109:25]
  wire [6:0] mmcm4_adv_DADDR; // @[Buf.scala 109:25]
  wire  mmcm4_adv_DEN; // @[Buf.scala 109:25]
  wire [15:0] mmcm4_adv_DI; // @[Buf.scala 109:25]
  wire  mmcm4_adv_DWE; // @[Buf.scala 109:25]
  wire  mmcm4_adv_PSCLK; // @[Buf.scala 109:25]
  wire  mmcm4_adv_PSEN; // @[Buf.scala 109:25]
  wire  mmcm4_adv_DCLK; // @[Buf.scala 109:25]
  wire  mmcm4_adv_PSINCDEC; // @[Buf.scala 109:25]
  wire  mmcm4_adv_LOCKED; // @[Buf.scala 109:25]
  wire  mmcm4_adv_CLKOUT0; // @[Buf.scala 109:25]
  wire  mmcm4_adv_CLKOUT1; // @[Buf.scala 109:25]
  wire  mmcm4_adv_CLKOUT2; // @[Buf.scala 109:25]
  wire  mmcm4_adv_CLKOUT3; // @[Buf.scala 109:25]
  wire  mmcm4_adv_CLKOUT4; // @[Buf.scala 109:25]
  wire  mmcm4_adv_CLKOUT5; // @[Buf.scala 109:25]
  wire  mmcm4_adv_CLKOUT6; // @[Buf.scala 109:25]
  MMCME4_ADV
    #(.CLKOUT5_DIVIDE(12.0), .CLKOUT3_DIVIDE(12.0), .CLKFBOUT_PHASE(0.0), .CLKIN1_PERIOD(10.0), .CLKOUT2_DIVIDE(12.0), .CLKOUT0_PHASE(0.0), .CLKFBOUT_MULT_F(12.0), .CLKOUT4_DIVIDE(12.0), .CLKOUT6_DIVIDE(2.0), .CLKOUT0_USE_FINE_PS("FALSE"), .COMPENSATION("INTERNAL"), .CLKOUT1_DIVIDE(12.0), .BANDWIDTH("OPTIMIZED"), .CLKFBOUT_USE_FINE_PS("FALSE"), .CLKOUT4_CASCADE("FALSE"), .CLKOUT0_DIVIDE_F(12.0), .CLKOUT0_DUTY_CYCLE(0.5), .REF_JITTER1(0.01), .DIVCLK_DIVIDE(1), .STARTUP_WAIT("FALSE"))
    mmcm4_adv ( // @[Buf.scala 109:25]
    .CLKIN1(mmcm4_adv_CLKIN1),
    .CLKIN2(mmcm4_adv_CLKIN2),
    .RST(mmcm4_adv_RST),
    .PWRDWN(mmcm4_adv_PWRDWN),
    .CDDCREQ(mmcm4_adv_CDDCREQ),
    .CLKINSEL(mmcm4_adv_CLKINSEL),
    .DADDR(mmcm4_adv_DADDR),
    .DEN(mmcm4_adv_DEN),
    .DI(mmcm4_adv_DI),
    .DWE(mmcm4_adv_DWE),
    .PSCLK(mmcm4_adv_PSCLK),
    .PSEN(mmcm4_adv_PSEN),
    .DCLK(mmcm4_adv_DCLK),
    .PSINCDEC(mmcm4_adv_PSINCDEC),
    .LOCKED(mmcm4_adv_LOCKED),
    .CLKOUT0(mmcm4_adv_CLKOUT0),
    .CLKOUT1(mmcm4_adv_CLKOUT1),
    .CLKOUT2(mmcm4_adv_CLKOUT2),
    .CLKOUT3(mmcm4_adv_CLKOUT3),
    .CLKOUT4(mmcm4_adv_CLKOUT4),
    .CLKOUT5(mmcm4_adv_CLKOUT5),
    .CLKOUT6(mmcm4_adv_CLKOUT6)
  );
  assign io_LOCKED = mmcm4_adv_LOCKED; // @[Buf.scala 123:25]
  assign io_CLKOUT0 = mmcm4_adv_CLKOUT0; // @[Buf.scala 124:26]
  assign io_CLKOUT1 = mmcm4_adv_CLKOUT1; // @[Buf.scala 125:26]
  assign io_CLKOUT2 = mmcm4_adv_CLKOUT2; // @[Buf.scala 126:26]
  assign io_CLKOUT3 = mmcm4_adv_CLKOUT3; // @[Buf.scala 127:26]
  assign io_CLKOUT4 = mmcm4_adv_CLKOUT4; // @[Buf.scala 128:26]
  assign io_CLKOUT5 = mmcm4_adv_CLKOUT5; // @[Buf.scala 129:26]
  assign mmcm4_adv_CLKIN1 = io_CLKIN1; // @[Buf.scala 121:25]
  assign mmcm4_adv_CLKIN2 = 1'h0; // @[Buf.scala 132:31]
  assign mmcm4_adv_RST = 1'h0; // @[Buf.scala 122:25]
  assign mmcm4_adv_PWRDWN = 1'h0; // @[Buf.scala 133:30]
  assign mmcm4_adv_CDDCREQ = 1'h0; // @[Buf.scala 134:32]
  assign mmcm4_adv_CLKINSEL = 1'h1; // @[Buf.scala 135:32]
  assign mmcm4_adv_DADDR = 7'h0; // @[Buf.scala 136:30]
  assign mmcm4_adv_DEN = 1'h0; // @[Buf.scala 137:28]
  assign mmcm4_adv_DI = 16'h0; // @[Buf.scala 138:26]
  assign mmcm4_adv_DWE = 1'h0; // @[Buf.scala 139:28]
  assign mmcm4_adv_PSCLK = 1'h0; // @[Buf.scala 140:30]
  assign mmcm4_adv_PSEN = 1'h0; // @[Buf.scala 141:28]
  assign mmcm4_adv_DCLK = 1'h0; // @[Buf.scala 142:28]
  assign mmcm4_adv_PSINCDEC = 1'h0; // @[Buf.scala 143:32]
endmodule
module MMCME4_ADV_Wrapper_1(
  input   io_CLKIN1,
  input   io_RST,
  output  io_LOCKED,
  output  io_CLKOUT0
);
  wire  mmcm4_adv_CLKIN1; // @[Buf.scala 109:25]
  wire  mmcm4_adv_CLKIN2; // @[Buf.scala 109:25]
  wire  mmcm4_adv_RST; // @[Buf.scala 109:25]
  wire  mmcm4_adv_PWRDWN; // @[Buf.scala 109:25]
  wire  mmcm4_adv_CDDCREQ; // @[Buf.scala 109:25]
  wire  mmcm4_adv_CLKINSEL; // @[Buf.scala 109:25]
  wire [6:0] mmcm4_adv_DADDR; // @[Buf.scala 109:25]
  wire  mmcm4_adv_DEN; // @[Buf.scala 109:25]
  wire [15:0] mmcm4_adv_DI; // @[Buf.scala 109:25]
  wire  mmcm4_adv_DWE; // @[Buf.scala 109:25]
  wire  mmcm4_adv_PSCLK; // @[Buf.scala 109:25]
  wire  mmcm4_adv_PSEN; // @[Buf.scala 109:25]
  wire  mmcm4_adv_DCLK; // @[Buf.scala 109:25]
  wire  mmcm4_adv_PSINCDEC; // @[Buf.scala 109:25]
  wire  mmcm4_adv_LOCKED; // @[Buf.scala 109:25]
  wire  mmcm4_adv_CLKOUT0; // @[Buf.scala 109:25]
  wire  mmcm4_adv_CLKOUT1; // @[Buf.scala 109:25]
  wire  mmcm4_adv_CLKOUT2; // @[Buf.scala 109:25]
  wire  mmcm4_adv_CLKOUT3; // @[Buf.scala 109:25]
  wire  mmcm4_adv_CLKOUT4; // @[Buf.scala 109:25]
  wire  mmcm4_adv_CLKOUT5; // @[Buf.scala 109:25]
  wire  mmcm4_adv_CLKOUT6; // @[Buf.scala 109:25]
  MMCME4_ADV
    #(.CLKOUT5_DIVIDE(2.0), .CLKOUT3_DIVIDE(2.0), .CLKFBOUT_PHASE(0.0), .CLKIN1_PERIOD(10.0), .CLKOUT2_DIVIDE(2.0), .CLKOUT0_PHASE(0.0), .CLKFBOUT_MULT_F(18.0), .CLKOUT4_DIVIDE(2.0), .CLKOUT6_DIVIDE(2.0), .CLKOUT0_USE_FINE_PS("FALSE"), .COMPENSATION("INTERNAL"), .CLKOUT1_DIVIDE(2.0), .BANDWIDTH("OPTIMIZED"), .CLKFBOUT_USE_FINE_PS("FALSE"), .CLKOUT4_CASCADE("FALSE"), .CLKOUT0_DIVIDE_F(2.0), .CLKOUT0_DUTY_CYCLE(0.5), .REF_JITTER1(0.01), .DIVCLK_DIVIDE(2), .STARTUP_WAIT("FALSE"))
    mmcm4_adv ( // @[Buf.scala 109:25]
    .CLKIN1(mmcm4_adv_CLKIN1),
    .CLKIN2(mmcm4_adv_CLKIN2),
    .RST(mmcm4_adv_RST),
    .PWRDWN(mmcm4_adv_PWRDWN),
    .CDDCREQ(mmcm4_adv_CDDCREQ),
    .CLKINSEL(mmcm4_adv_CLKINSEL),
    .DADDR(mmcm4_adv_DADDR),
    .DEN(mmcm4_adv_DEN),
    .DI(mmcm4_adv_DI),
    .DWE(mmcm4_adv_DWE),
    .PSCLK(mmcm4_adv_PSCLK),
    .PSEN(mmcm4_adv_PSEN),
    .DCLK(mmcm4_adv_DCLK),
    .PSINCDEC(mmcm4_adv_PSINCDEC),
    .LOCKED(mmcm4_adv_LOCKED),
    .CLKOUT0(mmcm4_adv_CLKOUT0),
    .CLKOUT1(mmcm4_adv_CLKOUT1),
    .CLKOUT2(mmcm4_adv_CLKOUT2),
    .CLKOUT3(mmcm4_adv_CLKOUT3),
    .CLKOUT4(mmcm4_adv_CLKOUT4),
    .CLKOUT5(mmcm4_adv_CLKOUT5),
    .CLKOUT6(mmcm4_adv_CLKOUT6)
  );
  assign io_LOCKED = mmcm4_adv_LOCKED; // @[Buf.scala 123:25]
  assign io_CLKOUT0 = mmcm4_adv_CLKOUT0; // @[Buf.scala 124:26]
  assign mmcm4_adv_CLKIN1 = io_CLKIN1; // @[Buf.scala 121:25]
  assign mmcm4_adv_CLKIN2 = 1'h0; // @[Buf.scala 132:31]
  assign mmcm4_adv_RST = io_RST; // @[Buf.scala 122:25]
  assign mmcm4_adv_PWRDWN = 1'h0; // @[Buf.scala 133:30]
  assign mmcm4_adv_CDDCREQ = 1'h0; // @[Buf.scala 134:32]
  assign mmcm4_adv_CLKINSEL = 1'h1; // @[Buf.scala 135:32]
  assign mmcm4_adv_DADDR = 7'h0; // @[Buf.scala 136:30]
  assign mmcm4_adv_DEN = 1'h0; // @[Buf.scala 137:28]
  assign mmcm4_adv_DI = 16'h0; // @[Buf.scala 138:26]
  assign mmcm4_adv_DWE = 1'h0; // @[Buf.scala 139:28]
  assign mmcm4_adv_PSCLK = 1'h0; // @[Buf.scala 140:30]
  assign mmcm4_adv_PSEN = 1'h0; // @[Buf.scala 141:28]
  assign mmcm4_adv_DCLK = 1'h0; // @[Buf.scala 142:28]
  assign mmcm4_adv_PSINCDEC = 1'h0; // @[Buf.scala 143:32]
endmodule
module HBM_DRIVER(
  input   clock,
  output  io_hbm_clk,
  output  io_hbm_rstn
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
`endif // RANDOMIZE_REG_INIT
  wire  mmcmGlbl_io_CLKIN1; // @[HBMDriver.scala 48:30]
  wire  mmcmGlbl_io_LOCKED; // @[HBMDriver.scala 48:30]
  wire  mmcmGlbl_io_CLKOUT0; // @[HBMDriver.scala 48:30]
  wire  mmcmGlbl_io_CLKOUT1; // @[HBMDriver.scala 48:30]
  wire  mmcmGlbl_io_CLKOUT2; // @[HBMDriver.scala 48:30]
  wire  mmcmGlbl_io_CLKOUT3; // @[HBMDriver.scala 48:30]
  wire  mmcmGlbl_io_CLKOUT4; // @[HBMDriver.scala 48:30]
  wire  mmcmGlbl_io_CLKOUT5; // @[HBMDriver.scala 48:30]
  wire  apb0Pclk_pad_O; // @[Buf.scala 33:34]
  wire  apb0Pclk_pad_I; // @[Buf.scala 33:34]
  wire  apb0Pclk_pad_1_O; // @[Buf.scala 17:34]
  wire  apb0Pclk_pad_1_I; // @[Buf.scala 17:34]
  wire  apb0Pclk_pad_2_O; // @[Buf.scala 33:34]
  wire  apb0Pclk_pad_2_I; // @[Buf.scala 33:34]
  wire  axiAclkIn0_pad_O; // @[Buf.scala 33:34]
  wire  axiAclkIn0_pad_I; // @[Buf.scala 33:34]
  wire  hbmRefClk0_pad_O; // @[Buf.scala 33:34]
  wire  hbmRefClk0_pad_I; // @[Buf.scala 33:34]
  wire  apb1Pclk_pad_O; // @[Buf.scala 33:34]
  wire  apb1Pclk_pad_I; // @[Buf.scala 33:34]
  wire  apb1Pclk_pad_1_O; // @[Buf.scala 17:34]
  wire  apb1Pclk_pad_1_I; // @[Buf.scala 17:34]
  wire  apb1Pclk_pad_2_O; // @[Buf.scala 33:34]
  wire  apb1Pclk_pad_2_I; // @[Buf.scala 33:34]
  wire  axiAclkIn1_pad_O; // @[Buf.scala 33:34]
  wire  axiAclkIn1_pad_I; // @[Buf.scala 33:34]
  wire  hbmRefClk1_pad_O; // @[Buf.scala 33:34]
  wire  hbmRefClk1_pad_I; // @[Buf.scala 33:34]
  wire  mmcmAxi_io_CLKIN1; // @[HBMDriver.scala 71:29]
  wire  mmcmAxi_io_RST; // @[HBMDriver.scala 71:29]
  wire  mmcmAxi_io_LOCKED; // @[HBMDriver.scala 71:29]
  wire  mmcmAxi_io_CLKOUT0; // @[HBMDriver.scala 71:29]
  wire  axiAclk_pad_O; // @[Buf.scala 33:34]
  wire  axiAclk_pad_I; // @[Buf.scala 33:34]
  wire  instHbm_HBM_REF_CLK_0; // @[HBMDriver.scala 92:29]
  wire  instHbm_HBM_REF_CLK_1; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_00_ACLK; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_00_ARESET_N; // @[HBMDriver.scala 92:29]
  wire [32:0] instHbm_AXI_00_ARADDR; // @[HBMDriver.scala 92:29]
  wire [1:0] instHbm_AXI_00_ARBURST; // @[HBMDriver.scala 92:29]
  wire [5:0] instHbm_AXI_00_ARID; // @[HBMDriver.scala 92:29]
  wire [3:0] instHbm_AXI_00_ARLEN; // @[HBMDriver.scala 92:29]
  wire [2:0] instHbm_AXI_00_ARSIZE; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_00_ARVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_00_ARREADY; // @[HBMDriver.scala 92:29]
  wire [32:0] instHbm_AXI_00_AWADDR; // @[HBMDriver.scala 92:29]
  wire [1:0] instHbm_AXI_00_AWBURST; // @[HBMDriver.scala 92:29]
  wire [5:0] instHbm_AXI_00_AWID; // @[HBMDriver.scala 92:29]
  wire [3:0] instHbm_AXI_00_AWLEN; // @[HBMDriver.scala 92:29]
  wire [2:0] instHbm_AXI_00_AWSIZE; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_00_AWVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_00_AWREADY; // @[HBMDriver.scala 92:29]
  wire [255:0] instHbm_AXI_00_WDATA; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_00_WLAST; // @[HBMDriver.scala 92:29]
  wire [31:0] instHbm_AXI_00_WSTRB; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_00_WVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_00_WREADY; // @[HBMDriver.scala 92:29]
  wire [255:0] instHbm_AXI_00_RDATA; // @[HBMDriver.scala 92:29]
  wire [5:0] instHbm_AXI_00_RID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_00_RLAST; // @[HBMDriver.scala 92:29]
  wire [1:0] instHbm_AXI_00_RRESP; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_00_RVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_00_RREADY; // @[HBMDriver.scala 92:29]
  wire [5:0] instHbm_AXI_00_BID; // @[HBMDriver.scala 92:29]
  wire [1:0] instHbm_AXI_00_BRESP; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_00_BVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_00_BREADY; // @[HBMDriver.scala 92:29]
  wire [31:0] instHbm_AXI_00_WDATA_PARITY; // @[HBMDriver.scala 92:29]
  wire [31:0] instHbm_AXI_00_RDATA_PARITY; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_01_ACLK; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_01_ARESET_N; // @[HBMDriver.scala 92:29]
  wire [32:0] instHbm_AXI_01_ARADDR; // @[HBMDriver.scala 92:29]
  wire [1:0] instHbm_AXI_01_ARBURST; // @[HBMDriver.scala 92:29]
  wire [5:0] instHbm_AXI_01_ARID; // @[HBMDriver.scala 92:29]
  wire [3:0] instHbm_AXI_01_ARLEN; // @[HBMDriver.scala 92:29]
  wire [2:0] instHbm_AXI_01_ARSIZE; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_01_ARVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_01_ARREADY; // @[HBMDriver.scala 92:29]
  wire [32:0] instHbm_AXI_01_AWADDR; // @[HBMDriver.scala 92:29]
  wire [1:0] instHbm_AXI_01_AWBURST; // @[HBMDriver.scala 92:29]
  wire [5:0] instHbm_AXI_01_AWID; // @[HBMDriver.scala 92:29]
  wire [3:0] instHbm_AXI_01_AWLEN; // @[HBMDriver.scala 92:29]
  wire [2:0] instHbm_AXI_01_AWSIZE; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_01_AWVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_01_AWREADY; // @[HBMDriver.scala 92:29]
  wire [255:0] instHbm_AXI_01_WDATA; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_01_WLAST; // @[HBMDriver.scala 92:29]
  wire [31:0] instHbm_AXI_01_WSTRB; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_01_WVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_01_WREADY; // @[HBMDriver.scala 92:29]
  wire [255:0] instHbm_AXI_01_RDATA; // @[HBMDriver.scala 92:29]
  wire [5:0] instHbm_AXI_01_RID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_01_RLAST; // @[HBMDriver.scala 92:29]
  wire [1:0] instHbm_AXI_01_RRESP; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_01_RVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_01_RREADY; // @[HBMDriver.scala 92:29]
  wire [5:0] instHbm_AXI_01_BID; // @[HBMDriver.scala 92:29]
  wire [1:0] instHbm_AXI_01_BRESP; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_01_BVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_01_BREADY; // @[HBMDriver.scala 92:29]
  wire [31:0] instHbm_AXI_01_WDATA_PARITY; // @[HBMDriver.scala 92:29]
  wire [31:0] instHbm_AXI_01_RDATA_PARITY; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_02_ACLK; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_02_ARESET_N; // @[HBMDriver.scala 92:29]
  wire [32:0] instHbm_AXI_02_ARADDR; // @[HBMDriver.scala 92:29]
  wire [1:0] instHbm_AXI_02_ARBURST; // @[HBMDriver.scala 92:29]
  wire [5:0] instHbm_AXI_02_ARID; // @[HBMDriver.scala 92:29]
  wire [3:0] instHbm_AXI_02_ARLEN; // @[HBMDriver.scala 92:29]
  wire [2:0] instHbm_AXI_02_ARSIZE; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_02_ARVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_02_ARREADY; // @[HBMDriver.scala 92:29]
  wire [32:0] instHbm_AXI_02_AWADDR; // @[HBMDriver.scala 92:29]
  wire [1:0] instHbm_AXI_02_AWBURST; // @[HBMDriver.scala 92:29]
  wire [5:0] instHbm_AXI_02_AWID; // @[HBMDriver.scala 92:29]
  wire [3:0] instHbm_AXI_02_AWLEN; // @[HBMDriver.scala 92:29]
  wire [2:0] instHbm_AXI_02_AWSIZE; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_02_AWVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_02_AWREADY; // @[HBMDriver.scala 92:29]
  wire [255:0] instHbm_AXI_02_WDATA; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_02_WLAST; // @[HBMDriver.scala 92:29]
  wire [31:0] instHbm_AXI_02_WSTRB; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_02_WVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_02_WREADY; // @[HBMDriver.scala 92:29]
  wire [255:0] instHbm_AXI_02_RDATA; // @[HBMDriver.scala 92:29]
  wire [5:0] instHbm_AXI_02_RID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_02_RLAST; // @[HBMDriver.scala 92:29]
  wire [1:0] instHbm_AXI_02_RRESP; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_02_RVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_02_RREADY; // @[HBMDriver.scala 92:29]
  wire [5:0] instHbm_AXI_02_BID; // @[HBMDriver.scala 92:29]
  wire [1:0] instHbm_AXI_02_BRESP; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_02_BVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_02_BREADY; // @[HBMDriver.scala 92:29]
  wire [31:0] instHbm_AXI_02_WDATA_PARITY; // @[HBMDriver.scala 92:29]
  wire [31:0] instHbm_AXI_02_RDATA_PARITY; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_03_ACLK; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_03_ARESET_N; // @[HBMDriver.scala 92:29]
  wire [32:0] instHbm_AXI_03_ARADDR; // @[HBMDriver.scala 92:29]
  wire [1:0] instHbm_AXI_03_ARBURST; // @[HBMDriver.scala 92:29]
  wire [5:0] instHbm_AXI_03_ARID; // @[HBMDriver.scala 92:29]
  wire [3:0] instHbm_AXI_03_ARLEN; // @[HBMDriver.scala 92:29]
  wire [2:0] instHbm_AXI_03_ARSIZE; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_03_ARVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_03_ARREADY; // @[HBMDriver.scala 92:29]
  wire [32:0] instHbm_AXI_03_AWADDR; // @[HBMDriver.scala 92:29]
  wire [1:0] instHbm_AXI_03_AWBURST; // @[HBMDriver.scala 92:29]
  wire [5:0] instHbm_AXI_03_AWID; // @[HBMDriver.scala 92:29]
  wire [3:0] instHbm_AXI_03_AWLEN; // @[HBMDriver.scala 92:29]
  wire [2:0] instHbm_AXI_03_AWSIZE; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_03_AWVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_03_AWREADY; // @[HBMDriver.scala 92:29]
  wire [255:0] instHbm_AXI_03_WDATA; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_03_WLAST; // @[HBMDriver.scala 92:29]
  wire [31:0] instHbm_AXI_03_WSTRB; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_03_WVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_03_WREADY; // @[HBMDriver.scala 92:29]
  wire [255:0] instHbm_AXI_03_RDATA; // @[HBMDriver.scala 92:29]
  wire [5:0] instHbm_AXI_03_RID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_03_RLAST; // @[HBMDriver.scala 92:29]
  wire [1:0] instHbm_AXI_03_RRESP; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_03_RVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_03_RREADY; // @[HBMDriver.scala 92:29]
  wire [5:0] instHbm_AXI_03_BID; // @[HBMDriver.scala 92:29]
  wire [1:0] instHbm_AXI_03_BRESP; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_03_BVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_03_BREADY; // @[HBMDriver.scala 92:29]
  wire [31:0] instHbm_AXI_03_WDATA_PARITY; // @[HBMDriver.scala 92:29]
  wire [31:0] instHbm_AXI_03_RDATA_PARITY; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_04_ACLK; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_04_ARESET_N; // @[HBMDriver.scala 92:29]
  wire [32:0] instHbm_AXI_04_ARADDR; // @[HBMDriver.scala 92:29]
  wire [1:0] instHbm_AXI_04_ARBURST; // @[HBMDriver.scala 92:29]
  wire [5:0] instHbm_AXI_04_ARID; // @[HBMDriver.scala 92:29]
  wire [3:0] instHbm_AXI_04_ARLEN; // @[HBMDriver.scala 92:29]
  wire [2:0] instHbm_AXI_04_ARSIZE; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_04_ARVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_04_ARREADY; // @[HBMDriver.scala 92:29]
  wire [32:0] instHbm_AXI_04_AWADDR; // @[HBMDriver.scala 92:29]
  wire [1:0] instHbm_AXI_04_AWBURST; // @[HBMDriver.scala 92:29]
  wire [5:0] instHbm_AXI_04_AWID; // @[HBMDriver.scala 92:29]
  wire [3:0] instHbm_AXI_04_AWLEN; // @[HBMDriver.scala 92:29]
  wire [2:0] instHbm_AXI_04_AWSIZE; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_04_AWVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_04_AWREADY; // @[HBMDriver.scala 92:29]
  wire [255:0] instHbm_AXI_04_WDATA; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_04_WLAST; // @[HBMDriver.scala 92:29]
  wire [31:0] instHbm_AXI_04_WSTRB; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_04_WVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_04_WREADY; // @[HBMDriver.scala 92:29]
  wire [255:0] instHbm_AXI_04_RDATA; // @[HBMDriver.scala 92:29]
  wire [5:0] instHbm_AXI_04_RID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_04_RLAST; // @[HBMDriver.scala 92:29]
  wire [1:0] instHbm_AXI_04_RRESP; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_04_RVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_04_RREADY; // @[HBMDriver.scala 92:29]
  wire [5:0] instHbm_AXI_04_BID; // @[HBMDriver.scala 92:29]
  wire [1:0] instHbm_AXI_04_BRESP; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_04_BVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_04_BREADY; // @[HBMDriver.scala 92:29]
  wire [31:0] instHbm_AXI_04_WDATA_PARITY; // @[HBMDriver.scala 92:29]
  wire [31:0] instHbm_AXI_04_RDATA_PARITY; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_05_ACLK; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_05_ARESET_N; // @[HBMDriver.scala 92:29]
  wire [32:0] instHbm_AXI_05_ARADDR; // @[HBMDriver.scala 92:29]
  wire [1:0] instHbm_AXI_05_ARBURST; // @[HBMDriver.scala 92:29]
  wire [5:0] instHbm_AXI_05_ARID; // @[HBMDriver.scala 92:29]
  wire [3:0] instHbm_AXI_05_ARLEN; // @[HBMDriver.scala 92:29]
  wire [2:0] instHbm_AXI_05_ARSIZE; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_05_ARVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_05_ARREADY; // @[HBMDriver.scala 92:29]
  wire [32:0] instHbm_AXI_05_AWADDR; // @[HBMDriver.scala 92:29]
  wire [1:0] instHbm_AXI_05_AWBURST; // @[HBMDriver.scala 92:29]
  wire [5:0] instHbm_AXI_05_AWID; // @[HBMDriver.scala 92:29]
  wire [3:0] instHbm_AXI_05_AWLEN; // @[HBMDriver.scala 92:29]
  wire [2:0] instHbm_AXI_05_AWSIZE; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_05_AWVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_05_AWREADY; // @[HBMDriver.scala 92:29]
  wire [255:0] instHbm_AXI_05_WDATA; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_05_WLAST; // @[HBMDriver.scala 92:29]
  wire [31:0] instHbm_AXI_05_WSTRB; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_05_WVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_05_WREADY; // @[HBMDriver.scala 92:29]
  wire [255:0] instHbm_AXI_05_RDATA; // @[HBMDriver.scala 92:29]
  wire [5:0] instHbm_AXI_05_RID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_05_RLAST; // @[HBMDriver.scala 92:29]
  wire [1:0] instHbm_AXI_05_RRESP; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_05_RVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_05_RREADY; // @[HBMDriver.scala 92:29]
  wire [5:0] instHbm_AXI_05_BID; // @[HBMDriver.scala 92:29]
  wire [1:0] instHbm_AXI_05_BRESP; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_05_BVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_05_BREADY; // @[HBMDriver.scala 92:29]
  wire [31:0] instHbm_AXI_05_WDATA_PARITY; // @[HBMDriver.scala 92:29]
  wire [31:0] instHbm_AXI_05_RDATA_PARITY; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_06_ACLK; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_06_ARESET_N; // @[HBMDriver.scala 92:29]
  wire [32:0] instHbm_AXI_06_ARADDR; // @[HBMDriver.scala 92:29]
  wire [1:0] instHbm_AXI_06_ARBURST; // @[HBMDriver.scala 92:29]
  wire [5:0] instHbm_AXI_06_ARID; // @[HBMDriver.scala 92:29]
  wire [3:0] instHbm_AXI_06_ARLEN; // @[HBMDriver.scala 92:29]
  wire [2:0] instHbm_AXI_06_ARSIZE; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_06_ARVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_06_ARREADY; // @[HBMDriver.scala 92:29]
  wire [32:0] instHbm_AXI_06_AWADDR; // @[HBMDriver.scala 92:29]
  wire [1:0] instHbm_AXI_06_AWBURST; // @[HBMDriver.scala 92:29]
  wire [5:0] instHbm_AXI_06_AWID; // @[HBMDriver.scala 92:29]
  wire [3:0] instHbm_AXI_06_AWLEN; // @[HBMDriver.scala 92:29]
  wire [2:0] instHbm_AXI_06_AWSIZE; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_06_AWVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_06_AWREADY; // @[HBMDriver.scala 92:29]
  wire [255:0] instHbm_AXI_06_WDATA; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_06_WLAST; // @[HBMDriver.scala 92:29]
  wire [31:0] instHbm_AXI_06_WSTRB; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_06_WVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_06_WREADY; // @[HBMDriver.scala 92:29]
  wire [255:0] instHbm_AXI_06_RDATA; // @[HBMDriver.scala 92:29]
  wire [5:0] instHbm_AXI_06_RID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_06_RLAST; // @[HBMDriver.scala 92:29]
  wire [1:0] instHbm_AXI_06_RRESP; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_06_RVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_06_RREADY; // @[HBMDriver.scala 92:29]
  wire [5:0] instHbm_AXI_06_BID; // @[HBMDriver.scala 92:29]
  wire [1:0] instHbm_AXI_06_BRESP; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_06_BVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_06_BREADY; // @[HBMDriver.scala 92:29]
  wire [31:0] instHbm_AXI_06_WDATA_PARITY; // @[HBMDriver.scala 92:29]
  wire [31:0] instHbm_AXI_06_RDATA_PARITY; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_07_ACLK; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_07_ARESET_N; // @[HBMDriver.scala 92:29]
  wire [32:0] instHbm_AXI_07_ARADDR; // @[HBMDriver.scala 92:29]
  wire [1:0] instHbm_AXI_07_ARBURST; // @[HBMDriver.scala 92:29]
  wire [5:0] instHbm_AXI_07_ARID; // @[HBMDriver.scala 92:29]
  wire [3:0] instHbm_AXI_07_ARLEN; // @[HBMDriver.scala 92:29]
  wire [2:0] instHbm_AXI_07_ARSIZE; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_07_ARVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_07_ARREADY; // @[HBMDriver.scala 92:29]
  wire [32:0] instHbm_AXI_07_AWADDR; // @[HBMDriver.scala 92:29]
  wire [1:0] instHbm_AXI_07_AWBURST; // @[HBMDriver.scala 92:29]
  wire [5:0] instHbm_AXI_07_AWID; // @[HBMDriver.scala 92:29]
  wire [3:0] instHbm_AXI_07_AWLEN; // @[HBMDriver.scala 92:29]
  wire [2:0] instHbm_AXI_07_AWSIZE; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_07_AWVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_07_AWREADY; // @[HBMDriver.scala 92:29]
  wire [255:0] instHbm_AXI_07_WDATA; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_07_WLAST; // @[HBMDriver.scala 92:29]
  wire [31:0] instHbm_AXI_07_WSTRB; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_07_WVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_07_WREADY; // @[HBMDriver.scala 92:29]
  wire [255:0] instHbm_AXI_07_RDATA; // @[HBMDriver.scala 92:29]
  wire [5:0] instHbm_AXI_07_RID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_07_RLAST; // @[HBMDriver.scala 92:29]
  wire [1:0] instHbm_AXI_07_RRESP; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_07_RVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_07_RREADY; // @[HBMDriver.scala 92:29]
  wire [5:0] instHbm_AXI_07_BID; // @[HBMDriver.scala 92:29]
  wire [1:0] instHbm_AXI_07_BRESP; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_07_BVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_07_BREADY; // @[HBMDriver.scala 92:29]
  wire [31:0] instHbm_AXI_07_WDATA_PARITY; // @[HBMDriver.scala 92:29]
  wire [31:0] instHbm_AXI_07_RDATA_PARITY; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_08_ACLK; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_08_ARESET_N; // @[HBMDriver.scala 92:29]
  wire [32:0] instHbm_AXI_08_ARADDR; // @[HBMDriver.scala 92:29]
  wire [1:0] instHbm_AXI_08_ARBURST; // @[HBMDriver.scala 92:29]
  wire [5:0] instHbm_AXI_08_ARID; // @[HBMDriver.scala 92:29]
  wire [3:0] instHbm_AXI_08_ARLEN; // @[HBMDriver.scala 92:29]
  wire [2:0] instHbm_AXI_08_ARSIZE; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_08_ARVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_08_ARREADY; // @[HBMDriver.scala 92:29]
  wire [32:0] instHbm_AXI_08_AWADDR; // @[HBMDriver.scala 92:29]
  wire [1:0] instHbm_AXI_08_AWBURST; // @[HBMDriver.scala 92:29]
  wire [5:0] instHbm_AXI_08_AWID; // @[HBMDriver.scala 92:29]
  wire [3:0] instHbm_AXI_08_AWLEN; // @[HBMDriver.scala 92:29]
  wire [2:0] instHbm_AXI_08_AWSIZE; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_08_AWVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_08_AWREADY; // @[HBMDriver.scala 92:29]
  wire [255:0] instHbm_AXI_08_WDATA; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_08_WLAST; // @[HBMDriver.scala 92:29]
  wire [31:0] instHbm_AXI_08_WSTRB; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_08_WVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_08_WREADY; // @[HBMDriver.scala 92:29]
  wire [255:0] instHbm_AXI_08_RDATA; // @[HBMDriver.scala 92:29]
  wire [5:0] instHbm_AXI_08_RID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_08_RLAST; // @[HBMDriver.scala 92:29]
  wire [1:0] instHbm_AXI_08_RRESP; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_08_RVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_08_RREADY; // @[HBMDriver.scala 92:29]
  wire [5:0] instHbm_AXI_08_BID; // @[HBMDriver.scala 92:29]
  wire [1:0] instHbm_AXI_08_BRESP; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_08_BVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_08_BREADY; // @[HBMDriver.scala 92:29]
  wire [31:0] instHbm_AXI_08_WDATA_PARITY; // @[HBMDriver.scala 92:29]
  wire [31:0] instHbm_AXI_08_RDATA_PARITY; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_09_ACLK; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_09_ARESET_N; // @[HBMDriver.scala 92:29]
  wire [32:0] instHbm_AXI_09_ARADDR; // @[HBMDriver.scala 92:29]
  wire [1:0] instHbm_AXI_09_ARBURST; // @[HBMDriver.scala 92:29]
  wire [5:0] instHbm_AXI_09_ARID; // @[HBMDriver.scala 92:29]
  wire [3:0] instHbm_AXI_09_ARLEN; // @[HBMDriver.scala 92:29]
  wire [2:0] instHbm_AXI_09_ARSIZE; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_09_ARVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_09_ARREADY; // @[HBMDriver.scala 92:29]
  wire [32:0] instHbm_AXI_09_AWADDR; // @[HBMDriver.scala 92:29]
  wire [1:0] instHbm_AXI_09_AWBURST; // @[HBMDriver.scala 92:29]
  wire [5:0] instHbm_AXI_09_AWID; // @[HBMDriver.scala 92:29]
  wire [3:0] instHbm_AXI_09_AWLEN; // @[HBMDriver.scala 92:29]
  wire [2:0] instHbm_AXI_09_AWSIZE; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_09_AWVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_09_AWREADY; // @[HBMDriver.scala 92:29]
  wire [255:0] instHbm_AXI_09_WDATA; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_09_WLAST; // @[HBMDriver.scala 92:29]
  wire [31:0] instHbm_AXI_09_WSTRB; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_09_WVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_09_WREADY; // @[HBMDriver.scala 92:29]
  wire [255:0] instHbm_AXI_09_RDATA; // @[HBMDriver.scala 92:29]
  wire [5:0] instHbm_AXI_09_RID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_09_RLAST; // @[HBMDriver.scala 92:29]
  wire [1:0] instHbm_AXI_09_RRESP; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_09_RVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_09_RREADY; // @[HBMDriver.scala 92:29]
  wire [5:0] instHbm_AXI_09_BID; // @[HBMDriver.scala 92:29]
  wire [1:0] instHbm_AXI_09_BRESP; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_09_BVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_09_BREADY; // @[HBMDriver.scala 92:29]
  wire [31:0] instHbm_AXI_09_WDATA_PARITY; // @[HBMDriver.scala 92:29]
  wire [31:0] instHbm_AXI_09_RDATA_PARITY; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_10_ACLK; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_10_ARESET_N; // @[HBMDriver.scala 92:29]
  wire [32:0] instHbm_AXI_10_ARADDR; // @[HBMDriver.scala 92:29]
  wire [1:0] instHbm_AXI_10_ARBURST; // @[HBMDriver.scala 92:29]
  wire [5:0] instHbm_AXI_10_ARID; // @[HBMDriver.scala 92:29]
  wire [3:0] instHbm_AXI_10_ARLEN; // @[HBMDriver.scala 92:29]
  wire [2:0] instHbm_AXI_10_ARSIZE; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_10_ARVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_10_ARREADY; // @[HBMDriver.scala 92:29]
  wire [32:0] instHbm_AXI_10_AWADDR; // @[HBMDriver.scala 92:29]
  wire [1:0] instHbm_AXI_10_AWBURST; // @[HBMDriver.scala 92:29]
  wire [5:0] instHbm_AXI_10_AWID; // @[HBMDriver.scala 92:29]
  wire [3:0] instHbm_AXI_10_AWLEN; // @[HBMDriver.scala 92:29]
  wire [2:0] instHbm_AXI_10_AWSIZE; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_10_AWVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_10_AWREADY; // @[HBMDriver.scala 92:29]
  wire [255:0] instHbm_AXI_10_WDATA; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_10_WLAST; // @[HBMDriver.scala 92:29]
  wire [31:0] instHbm_AXI_10_WSTRB; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_10_WVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_10_WREADY; // @[HBMDriver.scala 92:29]
  wire [255:0] instHbm_AXI_10_RDATA; // @[HBMDriver.scala 92:29]
  wire [5:0] instHbm_AXI_10_RID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_10_RLAST; // @[HBMDriver.scala 92:29]
  wire [1:0] instHbm_AXI_10_RRESP; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_10_RVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_10_RREADY; // @[HBMDriver.scala 92:29]
  wire [5:0] instHbm_AXI_10_BID; // @[HBMDriver.scala 92:29]
  wire [1:0] instHbm_AXI_10_BRESP; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_10_BVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_10_BREADY; // @[HBMDriver.scala 92:29]
  wire [31:0] instHbm_AXI_10_WDATA_PARITY; // @[HBMDriver.scala 92:29]
  wire [31:0] instHbm_AXI_10_RDATA_PARITY; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_11_ACLK; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_11_ARESET_N; // @[HBMDriver.scala 92:29]
  wire [32:0] instHbm_AXI_11_ARADDR; // @[HBMDriver.scala 92:29]
  wire [1:0] instHbm_AXI_11_ARBURST; // @[HBMDriver.scala 92:29]
  wire [5:0] instHbm_AXI_11_ARID; // @[HBMDriver.scala 92:29]
  wire [3:0] instHbm_AXI_11_ARLEN; // @[HBMDriver.scala 92:29]
  wire [2:0] instHbm_AXI_11_ARSIZE; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_11_ARVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_11_ARREADY; // @[HBMDriver.scala 92:29]
  wire [32:0] instHbm_AXI_11_AWADDR; // @[HBMDriver.scala 92:29]
  wire [1:0] instHbm_AXI_11_AWBURST; // @[HBMDriver.scala 92:29]
  wire [5:0] instHbm_AXI_11_AWID; // @[HBMDriver.scala 92:29]
  wire [3:0] instHbm_AXI_11_AWLEN; // @[HBMDriver.scala 92:29]
  wire [2:0] instHbm_AXI_11_AWSIZE; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_11_AWVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_11_AWREADY; // @[HBMDriver.scala 92:29]
  wire [255:0] instHbm_AXI_11_WDATA; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_11_WLAST; // @[HBMDriver.scala 92:29]
  wire [31:0] instHbm_AXI_11_WSTRB; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_11_WVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_11_WREADY; // @[HBMDriver.scala 92:29]
  wire [255:0] instHbm_AXI_11_RDATA; // @[HBMDriver.scala 92:29]
  wire [5:0] instHbm_AXI_11_RID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_11_RLAST; // @[HBMDriver.scala 92:29]
  wire [1:0] instHbm_AXI_11_RRESP; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_11_RVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_11_RREADY; // @[HBMDriver.scala 92:29]
  wire [5:0] instHbm_AXI_11_BID; // @[HBMDriver.scala 92:29]
  wire [1:0] instHbm_AXI_11_BRESP; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_11_BVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_11_BREADY; // @[HBMDriver.scala 92:29]
  wire [31:0] instHbm_AXI_11_WDATA_PARITY; // @[HBMDriver.scala 92:29]
  wire [31:0] instHbm_AXI_11_RDATA_PARITY; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_12_ACLK; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_12_ARESET_N; // @[HBMDriver.scala 92:29]
  wire [32:0] instHbm_AXI_12_ARADDR; // @[HBMDriver.scala 92:29]
  wire [1:0] instHbm_AXI_12_ARBURST; // @[HBMDriver.scala 92:29]
  wire [5:0] instHbm_AXI_12_ARID; // @[HBMDriver.scala 92:29]
  wire [3:0] instHbm_AXI_12_ARLEN; // @[HBMDriver.scala 92:29]
  wire [2:0] instHbm_AXI_12_ARSIZE; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_12_ARVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_12_ARREADY; // @[HBMDriver.scala 92:29]
  wire [32:0] instHbm_AXI_12_AWADDR; // @[HBMDriver.scala 92:29]
  wire [1:0] instHbm_AXI_12_AWBURST; // @[HBMDriver.scala 92:29]
  wire [5:0] instHbm_AXI_12_AWID; // @[HBMDriver.scala 92:29]
  wire [3:0] instHbm_AXI_12_AWLEN; // @[HBMDriver.scala 92:29]
  wire [2:0] instHbm_AXI_12_AWSIZE; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_12_AWVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_12_AWREADY; // @[HBMDriver.scala 92:29]
  wire [255:0] instHbm_AXI_12_WDATA; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_12_WLAST; // @[HBMDriver.scala 92:29]
  wire [31:0] instHbm_AXI_12_WSTRB; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_12_WVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_12_WREADY; // @[HBMDriver.scala 92:29]
  wire [255:0] instHbm_AXI_12_RDATA; // @[HBMDriver.scala 92:29]
  wire [5:0] instHbm_AXI_12_RID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_12_RLAST; // @[HBMDriver.scala 92:29]
  wire [1:0] instHbm_AXI_12_RRESP; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_12_RVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_12_RREADY; // @[HBMDriver.scala 92:29]
  wire [5:0] instHbm_AXI_12_BID; // @[HBMDriver.scala 92:29]
  wire [1:0] instHbm_AXI_12_BRESP; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_12_BVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_12_BREADY; // @[HBMDriver.scala 92:29]
  wire [31:0] instHbm_AXI_12_WDATA_PARITY; // @[HBMDriver.scala 92:29]
  wire [31:0] instHbm_AXI_12_RDATA_PARITY; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_13_ACLK; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_13_ARESET_N; // @[HBMDriver.scala 92:29]
  wire [32:0] instHbm_AXI_13_ARADDR; // @[HBMDriver.scala 92:29]
  wire [1:0] instHbm_AXI_13_ARBURST; // @[HBMDriver.scala 92:29]
  wire [5:0] instHbm_AXI_13_ARID; // @[HBMDriver.scala 92:29]
  wire [3:0] instHbm_AXI_13_ARLEN; // @[HBMDriver.scala 92:29]
  wire [2:0] instHbm_AXI_13_ARSIZE; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_13_ARVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_13_ARREADY; // @[HBMDriver.scala 92:29]
  wire [32:0] instHbm_AXI_13_AWADDR; // @[HBMDriver.scala 92:29]
  wire [1:0] instHbm_AXI_13_AWBURST; // @[HBMDriver.scala 92:29]
  wire [5:0] instHbm_AXI_13_AWID; // @[HBMDriver.scala 92:29]
  wire [3:0] instHbm_AXI_13_AWLEN; // @[HBMDriver.scala 92:29]
  wire [2:0] instHbm_AXI_13_AWSIZE; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_13_AWVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_13_AWREADY; // @[HBMDriver.scala 92:29]
  wire [255:0] instHbm_AXI_13_WDATA; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_13_WLAST; // @[HBMDriver.scala 92:29]
  wire [31:0] instHbm_AXI_13_WSTRB; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_13_WVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_13_WREADY; // @[HBMDriver.scala 92:29]
  wire [255:0] instHbm_AXI_13_RDATA; // @[HBMDriver.scala 92:29]
  wire [5:0] instHbm_AXI_13_RID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_13_RLAST; // @[HBMDriver.scala 92:29]
  wire [1:0] instHbm_AXI_13_RRESP; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_13_RVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_13_RREADY; // @[HBMDriver.scala 92:29]
  wire [5:0] instHbm_AXI_13_BID; // @[HBMDriver.scala 92:29]
  wire [1:0] instHbm_AXI_13_BRESP; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_13_BVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_13_BREADY; // @[HBMDriver.scala 92:29]
  wire [31:0] instHbm_AXI_13_WDATA_PARITY; // @[HBMDriver.scala 92:29]
  wire [31:0] instHbm_AXI_13_RDATA_PARITY; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_14_ACLK; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_14_ARESET_N; // @[HBMDriver.scala 92:29]
  wire [32:0] instHbm_AXI_14_ARADDR; // @[HBMDriver.scala 92:29]
  wire [1:0] instHbm_AXI_14_ARBURST; // @[HBMDriver.scala 92:29]
  wire [5:0] instHbm_AXI_14_ARID; // @[HBMDriver.scala 92:29]
  wire [3:0] instHbm_AXI_14_ARLEN; // @[HBMDriver.scala 92:29]
  wire [2:0] instHbm_AXI_14_ARSIZE; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_14_ARVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_14_ARREADY; // @[HBMDriver.scala 92:29]
  wire [32:0] instHbm_AXI_14_AWADDR; // @[HBMDriver.scala 92:29]
  wire [1:0] instHbm_AXI_14_AWBURST; // @[HBMDriver.scala 92:29]
  wire [5:0] instHbm_AXI_14_AWID; // @[HBMDriver.scala 92:29]
  wire [3:0] instHbm_AXI_14_AWLEN; // @[HBMDriver.scala 92:29]
  wire [2:0] instHbm_AXI_14_AWSIZE; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_14_AWVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_14_AWREADY; // @[HBMDriver.scala 92:29]
  wire [255:0] instHbm_AXI_14_WDATA; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_14_WLAST; // @[HBMDriver.scala 92:29]
  wire [31:0] instHbm_AXI_14_WSTRB; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_14_WVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_14_WREADY; // @[HBMDriver.scala 92:29]
  wire [255:0] instHbm_AXI_14_RDATA; // @[HBMDriver.scala 92:29]
  wire [5:0] instHbm_AXI_14_RID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_14_RLAST; // @[HBMDriver.scala 92:29]
  wire [1:0] instHbm_AXI_14_RRESP; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_14_RVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_14_RREADY; // @[HBMDriver.scala 92:29]
  wire [5:0] instHbm_AXI_14_BID; // @[HBMDriver.scala 92:29]
  wire [1:0] instHbm_AXI_14_BRESP; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_14_BVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_14_BREADY; // @[HBMDriver.scala 92:29]
  wire [31:0] instHbm_AXI_14_WDATA_PARITY; // @[HBMDriver.scala 92:29]
  wire [31:0] instHbm_AXI_14_RDATA_PARITY; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_15_ACLK; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_15_ARESET_N; // @[HBMDriver.scala 92:29]
  wire [32:0] instHbm_AXI_15_ARADDR; // @[HBMDriver.scala 92:29]
  wire [1:0] instHbm_AXI_15_ARBURST; // @[HBMDriver.scala 92:29]
  wire [5:0] instHbm_AXI_15_ARID; // @[HBMDriver.scala 92:29]
  wire [3:0] instHbm_AXI_15_ARLEN; // @[HBMDriver.scala 92:29]
  wire [2:0] instHbm_AXI_15_ARSIZE; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_15_ARVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_15_ARREADY; // @[HBMDriver.scala 92:29]
  wire [32:0] instHbm_AXI_15_AWADDR; // @[HBMDriver.scala 92:29]
  wire [1:0] instHbm_AXI_15_AWBURST; // @[HBMDriver.scala 92:29]
  wire [5:0] instHbm_AXI_15_AWID; // @[HBMDriver.scala 92:29]
  wire [3:0] instHbm_AXI_15_AWLEN; // @[HBMDriver.scala 92:29]
  wire [2:0] instHbm_AXI_15_AWSIZE; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_15_AWVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_15_AWREADY; // @[HBMDriver.scala 92:29]
  wire [255:0] instHbm_AXI_15_WDATA; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_15_WLAST; // @[HBMDriver.scala 92:29]
  wire [31:0] instHbm_AXI_15_WSTRB; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_15_WVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_15_WREADY; // @[HBMDriver.scala 92:29]
  wire [255:0] instHbm_AXI_15_RDATA; // @[HBMDriver.scala 92:29]
  wire [5:0] instHbm_AXI_15_RID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_15_RLAST; // @[HBMDriver.scala 92:29]
  wire [1:0] instHbm_AXI_15_RRESP; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_15_RVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_15_RREADY; // @[HBMDriver.scala 92:29]
  wire [5:0] instHbm_AXI_15_BID; // @[HBMDriver.scala 92:29]
  wire [1:0] instHbm_AXI_15_BRESP; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_15_BVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_15_BREADY; // @[HBMDriver.scala 92:29]
  wire [31:0] instHbm_AXI_15_WDATA_PARITY; // @[HBMDriver.scala 92:29]
  wire [31:0] instHbm_AXI_15_RDATA_PARITY; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_16_ACLK; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_16_ARESET_N; // @[HBMDriver.scala 92:29]
  wire [32:0] instHbm_AXI_16_ARADDR; // @[HBMDriver.scala 92:29]
  wire [1:0] instHbm_AXI_16_ARBURST; // @[HBMDriver.scala 92:29]
  wire [5:0] instHbm_AXI_16_ARID; // @[HBMDriver.scala 92:29]
  wire [3:0] instHbm_AXI_16_ARLEN; // @[HBMDriver.scala 92:29]
  wire [2:0] instHbm_AXI_16_ARSIZE; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_16_ARVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_16_ARREADY; // @[HBMDriver.scala 92:29]
  wire [32:0] instHbm_AXI_16_AWADDR; // @[HBMDriver.scala 92:29]
  wire [1:0] instHbm_AXI_16_AWBURST; // @[HBMDriver.scala 92:29]
  wire [5:0] instHbm_AXI_16_AWID; // @[HBMDriver.scala 92:29]
  wire [3:0] instHbm_AXI_16_AWLEN; // @[HBMDriver.scala 92:29]
  wire [2:0] instHbm_AXI_16_AWSIZE; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_16_AWVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_16_AWREADY; // @[HBMDriver.scala 92:29]
  wire [255:0] instHbm_AXI_16_WDATA; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_16_WLAST; // @[HBMDriver.scala 92:29]
  wire [31:0] instHbm_AXI_16_WSTRB; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_16_WVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_16_WREADY; // @[HBMDriver.scala 92:29]
  wire [255:0] instHbm_AXI_16_RDATA; // @[HBMDriver.scala 92:29]
  wire [5:0] instHbm_AXI_16_RID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_16_RLAST; // @[HBMDriver.scala 92:29]
  wire [1:0] instHbm_AXI_16_RRESP; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_16_RVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_16_RREADY; // @[HBMDriver.scala 92:29]
  wire [5:0] instHbm_AXI_16_BID; // @[HBMDriver.scala 92:29]
  wire [1:0] instHbm_AXI_16_BRESP; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_16_BVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_16_BREADY; // @[HBMDriver.scala 92:29]
  wire [31:0] instHbm_AXI_16_WDATA_PARITY; // @[HBMDriver.scala 92:29]
  wire [31:0] instHbm_AXI_16_RDATA_PARITY; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_17_ACLK; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_17_ARESET_N; // @[HBMDriver.scala 92:29]
  wire [32:0] instHbm_AXI_17_ARADDR; // @[HBMDriver.scala 92:29]
  wire [1:0] instHbm_AXI_17_ARBURST; // @[HBMDriver.scala 92:29]
  wire [5:0] instHbm_AXI_17_ARID; // @[HBMDriver.scala 92:29]
  wire [3:0] instHbm_AXI_17_ARLEN; // @[HBMDriver.scala 92:29]
  wire [2:0] instHbm_AXI_17_ARSIZE; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_17_ARVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_17_ARREADY; // @[HBMDriver.scala 92:29]
  wire [32:0] instHbm_AXI_17_AWADDR; // @[HBMDriver.scala 92:29]
  wire [1:0] instHbm_AXI_17_AWBURST; // @[HBMDriver.scala 92:29]
  wire [5:0] instHbm_AXI_17_AWID; // @[HBMDriver.scala 92:29]
  wire [3:0] instHbm_AXI_17_AWLEN; // @[HBMDriver.scala 92:29]
  wire [2:0] instHbm_AXI_17_AWSIZE; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_17_AWVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_17_AWREADY; // @[HBMDriver.scala 92:29]
  wire [255:0] instHbm_AXI_17_WDATA; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_17_WLAST; // @[HBMDriver.scala 92:29]
  wire [31:0] instHbm_AXI_17_WSTRB; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_17_WVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_17_WREADY; // @[HBMDriver.scala 92:29]
  wire [255:0] instHbm_AXI_17_RDATA; // @[HBMDriver.scala 92:29]
  wire [5:0] instHbm_AXI_17_RID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_17_RLAST; // @[HBMDriver.scala 92:29]
  wire [1:0] instHbm_AXI_17_RRESP; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_17_RVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_17_RREADY; // @[HBMDriver.scala 92:29]
  wire [5:0] instHbm_AXI_17_BID; // @[HBMDriver.scala 92:29]
  wire [1:0] instHbm_AXI_17_BRESP; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_17_BVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_17_BREADY; // @[HBMDriver.scala 92:29]
  wire [31:0] instHbm_AXI_17_WDATA_PARITY; // @[HBMDriver.scala 92:29]
  wire [31:0] instHbm_AXI_17_RDATA_PARITY; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_18_ACLK; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_18_ARESET_N; // @[HBMDriver.scala 92:29]
  wire [32:0] instHbm_AXI_18_ARADDR; // @[HBMDriver.scala 92:29]
  wire [1:0] instHbm_AXI_18_ARBURST; // @[HBMDriver.scala 92:29]
  wire [5:0] instHbm_AXI_18_ARID; // @[HBMDriver.scala 92:29]
  wire [3:0] instHbm_AXI_18_ARLEN; // @[HBMDriver.scala 92:29]
  wire [2:0] instHbm_AXI_18_ARSIZE; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_18_ARVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_18_ARREADY; // @[HBMDriver.scala 92:29]
  wire [32:0] instHbm_AXI_18_AWADDR; // @[HBMDriver.scala 92:29]
  wire [1:0] instHbm_AXI_18_AWBURST; // @[HBMDriver.scala 92:29]
  wire [5:0] instHbm_AXI_18_AWID; // @[HBMDriver.scala 92:29]
  wire [3:0] instHbm_AXI_18_AWLEN; // @[HBMDriver.scala 92:29]
  wire [2:0] instHbm_AXI_18_AWSIZE; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_18_AWVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_18_AWREADY; // @[HBMDriver.scala 92:29]
  wire [255:0] instHbm_AXI_18_WDATA; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_18_WLAST; // @[HBMDriver.scala 92:29]
  wire [31:0] instHbm_AXI_18_WSTRB; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_18_WVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_18_WREADY; // @[HBMDriver.scala 92:29]
  wire [255:0] instHbm_AXI_18_RDATA; // @[HBMDriver.scala 92:29]
  wire [5:0] instHbm_AXI_18_RID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_18_RLAST; // @[HBMDriver.scala 92:29]
  wire [1:0] instHbm_AXI_18_RRESP; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_18_RVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_18_RREADY; // @[HBMDriver.scala 92:29]
  wire [5:0] instHbm_AXI_18_BID; // @[HBMDriver.scala 92:29]
  wire [1:0] instHbm_AXI_18_BRESP; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_18_BVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_18_BREADY; // @[HBMDriver.scala 92:29]
  wire [31:0] instHbm_AXI_18_WDATA_PARITY; // @[HBMDriver.scala 92:29]
  wire [31:0] instHbm_AXI_18_RDATA_PARITY; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_19_ACLK; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_19_ARESET_N; // @[HBMDriver.scala 92:29]
  wire [32:0] instHbm_AXI_19_ARADDR; // @[HBMDriver.scala 92:29]
  wire [1:0] instHbm_AXI_19_ARBURST; // @[HBMDriver.scala 92:29]
  wire [5:0] instHbm_AXI_19_ARID; // @[HBMDriver.scala 92:29]
  wire [3:0] instHbm_AXI_19_ARLEN; // @[HBMDriver.scala 92:29]
  wire [2:0] instHbm_AXI_19_ARSIZE; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_19_ARVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_19_ARREADY; // @[HBMDriver.scala 92:29]
  wire [32:0] instHbm_AXI_19_AWADDR; // @[HBMDriver.scala 92:29]
  wire [1:0] instHbm_AXI_19_AWBURST; // @[HBMDriver.scala 92:29]
  wire [5:0] instHbm_AXI_19_AWID; // @[HBMDriver.scala 92:29]
  wire [3:0] instHbm_AXI_19_AWLEN; // @[HBMDriver.scala 92:29]
  wire [2:0] instHbm_AXI_19_AWSIZE; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_19_AWVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_19_AWREADY; // @[HBMDriver.scala 92:29]
  wire [255:0] instHbm_AXI_19_WDATA; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_19_WLAST; // @[HBMDriver.scala 92:29]
  wire [31:0] instHbm_AXI_19_WSTRB; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_19_WVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_19_WREADY; // @[HBMDriver.scala 92:29]
  wire [255:0] instHbm_AXI_19_RDATA; // @[HBMDriver.scala 92:29]
  wire [5:0] instHbm_AXI_19_RID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_19_RLAST; // @[HBMDriver.scala 92:29]
  wire [1:0] instHbm_AXI_19_RRESP; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_19_RVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_19_RREADY; // @[HBMDriver.scala 92:29]
  wire [5:0] instHbm_AXI_19_BID; // @[HBMDriver.scala 92:29]
  wire [1:0] instHbm_AXI_19_BRESP; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_19_BVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_19_BREADY; // @[HBMDriver.scala 92:29]
  wire [31:0] instHbm_AXI_19_WDATA_PARITY; // @[HBMDriver.scala 92:29]
  wire [31:0] instHbm_AXI_19_RDATA_PARITY; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_20_ACLK; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_20_ARESET_N; // @[HBMDriver.scala 92:29]
  wire [32:0] instHbm_AXI_20_ARADDR; // @[HBMDriver.scala 92:29]
  wire [1:0] instHbm_AXI_20_ARBURST; // @[HBMDriver.scala 92:29]
  wire [5:0] instHbm_AXI_20_ARID; // @[HBMDriver.scala 92:29]
  wire [3:0] instHbm_AXI_20_ARLEN; // @[HBMDriver.scala 92:29]
  wire [2:0] instHbm_AXI_20_ARSIZE; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_20_ARVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_20_ARREADY; // @[HBMDriver.scala 92:29]
  wire [32:0] instHbm_AXI_20_AWADDR; // @[HBMDriver.scala 92:29]
  wire [1:0] instHbm_AXI_20_AWBURST; // @[HBMDriver.scala 92:29]
  wire [5:0] instHbm_AXI_20_AWID; // @[HBMDriver.scala 92:29]
  wire [3:0] instHbm_AXI_20_AWLEN; // @[HBMDriver.scala 92:29]
  wire [2:0] instHbm_AXI_20_AWSIZE; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_20_AWVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_20_AWREADY; // @[HBMDriver.scala 92:29]
  wire [255:0] instHbm_AXI_20_WDATA; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_20_WLAST; // @[HBMDriver.scala 92:29]
  wire [31:0] instHbm_AXI_20_WSTRB; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_20_WVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_20_WREADY; // @[HBMDriver.scala 92:29]
  wire [255:0] instHbm_AXI_20_RDATA; // @[HBMDriver.scala 92:29]
  wire [5:0] instHbm_AXI_20_RID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_20_RLAST; // @[HBMDriver.scala 92:29]
  wire [1:0] instHbm_AXI_20_RRESP; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_20_RVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_20_RREADY; // @[HBMDriver.scala 92:29]
  wire [5:0] instHbm_AXI_20_BID; // @[HBMDriver.scala 92:29]
  wire [1:0] instHbm_AXI_20_BRESP; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_20_BVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_20_BREADY; // @[HBMDriver.scala 92:29]
  wire [31:0] instHbm_AXI_20_WDATA_PARITY; // @[HBMDriver.scala 92:29]
  wire [31:0] instHbm_AXI_20_RDATA_PARITY; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_21_ACLK; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_21_ARESET_N; // @[HBMDriver.scala 92:29]
  wire [32:0] instHbm_AXI_21_ARADDR; // @[HBMDriver.scala 92:29]
  wire [1:0] instHbm_AXI_21_ARBURST; // @[HBMDriver.scala 92:29]
  wire [5:0] instHbm_AXI_21_ARID; // @[HBMDriver.scala 92:29]
  wire [3:0] instHbm_AXI_21_ARLEN; // @[HBMDriver.scala 92:29]
  wire [2:0] instHbm_AXI_21_ARSIZE; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_21_ARVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_21_ARREADY; // @[HBMDriver.scala 92:29]
  wire [32:0] instHbm_AXI_21_AWADDR; // @[HBMDriver.scala 92:29]
  wire [1:0] instHbm_AXI_21_AWBURST; // @[HBMDriver.scala 92:29]
  wire [5:0] instHbm_AXI_21_AWID; // @[HBMDriver.scala 92:29]
  wire [3:0] instHbm_AXI_21_AWLEN; // @[HBMDriver.scala 92:29]
  wire [2:0] instHbm_AXI_21_AWSIZE; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_21_AWVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_21_AWREADY; // @[HBMDriver.scala 92:29]
  wire [255:0] instHbm_AXI_21_WDATA; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_21_WLAST; // @[HBMDriver.scala 92:29]
  wire [31:0] instHbm_AXI_21_WSTRB; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_21_WVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_21_WREADY; // @[HBMDriver.scala 92:29]
  wire [255:0] instHbm_AXI_21_RDATA; // @[HBMDriver.scala 92:29]
  wire [5:0] instHbm_AXI_21_RID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_21_RLAST; // @[HBMDriver.scala 92:29]
  wire [1:0] instHbm_AXI_21_RRESP; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_21_RVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_21_RREADY; // @[HBMDriver.scala 92:29]
  wire [5:0] instHbm_AXI_21_BID; // @[HBMDriver.scala 92:29]
  wire [1:0] instHbm_AXI_21_BRESP; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_21_BVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_21_BREADY; // @[HBMDriver.scala 92:29]
  wire [31:0] instHbm_AXI_21_WDATA_PARITY; // @[HBMDriver.scala 92:29]
  wire [31:0] instHbm_AXI_21_RDATA_PARITY; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_22_ACLK; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_22_ARESET_N; // @[HBMDriver.scala 92:29]
  wire [32:0] instHbm_AXI_22_ARADDR; // @[HBMDriver.scala 92:29]
  wire [1:0] instHbm_AXI_22_ARBURST; // @[HBMDriver.scala 92:29]
  wire [5:0] instHbm_AXI_22_ARID; // @[HBMDriver.scala 92:29]
  wire [3:0] instHbm_AXI_22_ARLEN; // @[HBMDriver.scala 92:29]
  wire [2:0] instHbm_AXI_22_ARSIZE; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_22_ARVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_22_ARREADY; // @[HBMDriver.scala 92:29]
  wire [32:0] instHbm_AXI_22_AWADDR; // @[HBMDriver.scala 92:29]
  wire [1:0] instHbm_AXI_22_AWBURST; // @[HBMDriver.scala 92:29]
  wire [5:0] instHbm_AXI_22_AWID; // @[HBMDriver.scala 92:29]
  wire [3:0] instHbm_AXI_22_AWLEN; // @[HBMDriver.scala 92:29]
  wire [2:0] instHbm_AXI_22_AWSIZE; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_22_AWVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_22_AWREADY; // @[HBMDriver.scala 92:29]
  wire [255:0] instHbm_AXI_22_WDATA; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_22_WLAST; // @[HBMDriver.scala 92:29]
  wire [31:0] instHbm_AXI_22_WSTRB; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_22_WVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_22_WREADY; // @[HBMDriver.scala 92:29]
  wire [255:0] instHbm_AXI_22_RDATA; // @[HBMDriver.scala 92:29]
  wire [5:0] instHbm_AXI_22_RID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_22_RLAST; // @[HBMDriver.scala 92:29]
  wire [1:0] instHbm_AXI_22_RRESP; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_22_RVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_22_RREADY; // @[HBMDriver.scala 92:29]
  wire [5:0] instHbm_AXI_22_BID; // @[HBMDriver.scala 92:29]
  wire [1:0] instHbm_AXI_22_BRESP; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_22_BVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_22_BREADY; // @[HBMDriver.scala 92:29]
  wire [31:0] instHbm_AXI_22_WDATA_PARITY; // @[HBMDriver.scala 92:29]
  wire [31:0] instHbm_AXI_22_RDATA_PARITY; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_23_ACLK; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_23_ARESET_N; // @[HBMDriver.scala 92:29]
  wire [32:0] instHbm_AXI_23_ARADDR; // @[HBMDriver.scala 92:29]
  wire [1:0] instHbm_AXI_23_ARBURST; // @[HBMDriver.scala 92:29]
  wire [5:0] instHbm_AXI_23_ARID; // @[HBMDriver.scala 92:29]
  wire [3:0] instHbm_AXI_23_ARLEN; // @[HBMDriver.scala 92:29]
  wire [2:0] instHbm_AXI_23_ARSIZE; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_23_ARVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_23_ARREADY; // @[HBMDriver.scala 92:29]
  wire [32:0] instHbm_AXI_23_AWADDR; // @[HBMDriver.scala 92:29]
  wire [1:0] instHbm_AXI_23_AWBURST; // @[HBMDriver.scala 92:29]
  wire [5:0] instHbm_AXI_23_AWID; // @[HBMDriver.scala 92:29]
  wire [3:0] instHbm_AXI_23_AWLEN; // @[HBMDriver.scala 92:29]
  wire [2:0] instHbm_AXI_23_AWSIZE; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_23_AWVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_23_AWREADY; // @[HBMDriver.scala 92:29]
  wire [255:0] instHbm_AXI_23_WDATA; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_23_WLAST; // @[HBMDriver.scala 92:29]
  wire [31:0] instHbm_AXI_23_WSTRB; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_23_WVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_23_WREADY; // @[HBMDriver.scala 92:29]
  wire [255:0] instHbm_AXI_23_RDATA; // @[HBMDriver.scala 92:29]
  wire [5:0] instHbm_AXI_23_RID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_23_RLAST; // @[HBMDriver.scala 92:29]
  wire [1:0] instHbm_AXI_23_RRESP; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_23_RVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_23_RREADY; // @[HBMDriver.scala 92:29]
  wire [5:0] instHbm_AXI_23_BID; // @[HBMDriver.scala 92:29]
  wire [1:0] instHbm_AXI_23_BRESP; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_23_BVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_23_BREADY; // @[HBMDriver.scala 92:29]
  wire [31:0] instHbm_AXI_23_WDATA_PARITY; // @[HBMDriver.scala 92:29]
  wire [31:0] instHbm_AXI_23_RDATA_PARITY; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_24_ACLK; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_24_ARESET_N; // @[HBMDriver.scala 92:29]
  wire [32:0] instHbm_AXI_24_ARADDR; // @[HBMDriver.scala 92:29]
  wire [1:0] instHbm_AXI_24_ARBURST; // @[HBMDriver.scala 92:29]
  wire [5:0] instHbm_AXI_24_ARID; // @[HBMDriver.scala 92:29]
  wire [3:0] instHbm_AXI_24_ARLEN; // @[HBMDriver.scala 92:29]
  wire [2:0] instHbm_AXI_24_ARSIZE; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_24_ARVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_24_ARREADY; // @[HBMDriver.scala 92:29]
  wire [32:0] instHbm_AXI_24_AWADDR; // @[HBMDriver.scala 92:29]
  wire [1:0] instHbm_AXI_24_AWBURST; // @[HBMDriver.scala 92:29]
  wire [5:0] instHbm_AXI_24_AWID; // @[HBMDriver.scala 92:29]
  wire [3:0] instHbm_AXI_24_AWLEN; // @[HBMDriver.scala 92:29]
  wire [2:0] instHbm_AXI_24_AWSIZE; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_24_AWVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_24_AWREADY; // @[HBMDriver.scala 92:29]
  wire [255:0] instHbm_AXI_24_WDATA; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_24_WLAST; // @[HBMDriver.scala 92:29]
  wire [31:0] instHbm_AXI_24_WSTRB; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_24_WVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_24_WREADY; // @[HBMDriver.scala 92:29]
  wire [255:0] instHbm_AXI_24_RDATA; // @[HBMDriver.scala 92:29]
  wire [5:0] instHbm_AXI_24_RID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_24_RLAST; // @[HBMDriver.scala 92:29]
  wire [1:0] instHbm_AXI_24_RRESP; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_24_RVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_24_RREADY; // @[HBMDriver.scala 92:29]
  wire [5:0] instHbm_AXI_24_BID; // @[HBMDriver.scala 92:29]
  wire [1:0] instHbm_AXI_24_BRESP; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_24_BVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_24_BREADY; // @[HBMDriver.scala 92:29]
  wire [31:0] instHbm_AXI_24_WDATA_PARITY; // @[HBMDriver.scala 92:29]
  wire [31:0] instHbm_AXI_24_RDATA_PARITY; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_25_ACLK; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_25_ARESET_N; // @[HBMDriver.scala 92:29]
  wire [32:0] instHbm_AXI_25_ARADDR; // @[HBMDriver.scala 92:29]
  wire [1:0] instHbm_AXI_25_ARBURST; // @[HBMDriver.scala 92:29]
  wire [5:0] instHbm_AXI_25_ARID; // @[HBMDriver.scala 92:29]
  wire [3:0] instHbm_AXI_25_ARLEN; // @[HBMDriver.scala 92:29]
  wire [2:0] instHbm_AXI_25_ARSIZE; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_25_ARVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_25_ARREADY; // @[HBMDriver.scala 92:29]
  wire [32:0] instHbm_AXI_25_AWADDR; // @[HBMDriver.scala 92:29]
  wire [1:0] instHbm_AXI_25_AWBURST; // @[HBMDriver.scala 92:29]
  wire [5:0] instHbm_AXI_25_AWID; // @[HBMDriver.scala 92:29]
  wire [3:0] instHbm_AXI_25_AWLEN; // @[HBMDriver.scala 92:29]
  wire [2:0] instHbm_AXI_25_AWSIZE; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_25_AWVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_25_AWREADY; // @[HBMDriver.scala 92:29]
  wire [255:0] instHbm_AXI_25_WDATA; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_25_WLAST; // @[HBMDriver.scala 92:29]
  wire [31:0] instHbm_AXI_25_WSTRB; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_25_WVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_25_WREADY; // @[HBMDriver.scala 92:29]
  wire [255:0] instHbm_AXI_25_RDATA; // @[HBMDriver.scala 92:29]
  wire [5:0] instHbm_AXI_25_RID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_25_RLAST; // @[HBMDriver.scala 92:29]
  wire [1:0] instHbm_AXI_25_RRESP; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_25_RVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_25_RREADY; // @[HBMDriver.scala 92:29]
  wire [5:0] instHbm_AXI_25_BID; // @[HBMDriver.scala 92:29]
  wire [1:0] instHbm_AXI_25_BRESP; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_25_BVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_25_BREADY; // @[HBMDriver.scala 92:29]
  wire [31:0] instHbm_AXI_25_WDATA_PARITY; // @[HBMDriver.scala 92:29]
  wire [31:0] instHbm_AXI_25_RDATA_PARITY; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_26_ACLK; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_26_ARESET_N; // @[HBMDriver.scala 92:29]
  wire [32:0] instHbm_AXI_26_ARADDR; // @[HBMDriver.scala 92:29]
  wire [1:0] instHbm_AXI_26_ARBURST; // @[HBMDriver.scala 92:29]
  wire [5:0] instHbm_AXI_26_ARID; // @[HBMDriver.scala 92:29]
  wire [3:0] instHbm_AXI_26_ARLEN; // @[HBMDriver.scala 92:29]
  wire [2:0] instHbm_AXI_26_ARSIZE; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_26_ARVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_26_ARREADY; // @[HBMDriver.scala 92:29]
  wire [32:0] instHbm_AXI_26_AWADDR; // @[HBMDriver.scala 92:29]
  wire [1:0] instHbm_AXI_26_AWBURST; // @[HBMDriver.scala 92:29]
  wire [5:0] instHbm_AXI_26_AWID; // @[HBMDriver.scala 92:29]
  wire [3:0] instHbm_AXI_26_AWLEN; // @[HBMDriver.scala 92:29]
  wire [2:0] instHbm_AXI_26_AWSIZE; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_26_AWVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_26_AWREADY; // @[HBMDriver.scala 92:29]
  wire [255:0] instHbm_AXI_26_WDATA; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_26_WLAST; // @[HBMDriver.scala 92:29]
  wire [31:0] instHbm_AXI_26_WSTRB; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_26_WVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_26_WREADY; // @[HBMDriver.scala 92:29]
  wire [255:0] instHbm_AXI_26_RDATA; // @[HBMDriver.scala 92:29]
  wire [5:0] instHbm_AXI_26_RID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_26_RLAST; // @[HBMDriver.scala 92:29]
  wire [1:0] instHbm_AXI_26_RRESP; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_26_RVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_26_RREADY; // @[HBMDriver.scala 92:29]
  wire [5:0] instHbm_AXI_26_BID; // @[HBMDriver.scala 92:29]
  wire [1:0] instHbm_AXI_26_BRESP; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_26_BVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_26_BREADY; // @[HBMDriver.scala 92:29]
  wire [31:0] instHbm_AXI_26_WDATA_PARITY; // @[HBMDriver.scala 92:29]
  wire [31:0] instHbm_AXI_26_RDATA_PARITY; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_27_ACLK; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_27_ARESET_N; // @[HBMDriver.scala 92:29]
  wire [32:0] instHbm_AXI_27_ARADDR; // @[HBMDriver.scala 92:29]
  wire [1:0] instHbm_AXI_27_ARBURST; // @[HBMDriver.scala 92:29]
  wire [5:0] instHbm_AXI_27_ARID; // @[HBMDriver.scala 92:29]
  wire [3:0] instHbm_AXI_27_ARLEN; // @[HBMDriver.scala 92:29]
  wire [2:0] instHbm_AXI_27_ARSIZE; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_27_ARVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_27_ARREADY; // @[HBMDriver.scala 92:29]
  wire [32:0] instHbm_AXI_27_AWADDR; // @[HBMDriver.scala 92:29]
  wire [1:0] instHbm_AXI_27_AWBURST; // @[HBMDriver.scala 92:29]
  wire [5:0] instHbm_AXI_27_AWID; // @[HBMDriver.scala 92:29]
  wire [3:0] instHbm_AXI_27_AWLEN; // @[HBMDriver.scala 92:29]
  wire [2:0] instHbm_AXI_27_AWSIZE; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_27_AWVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_27_AWREADY; // @[HBMDriver.scala 92:29]
  wire [255:0] instHbm_AXI_27_WDATA; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_27_WLAST; // @[HBMDriver.scala 92:29]
  wire [31:0] instHbm_AXI_27_WSTRB; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_27_WVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_27_WREADY; // @[HBMDriver.scala 92:29]
  wire [255:0] instHbm_AXI_27_RDATA; // @[HBMDriver.scala 92:29]
  wire [5:0] instHbm_AXI_27_RID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_27_RLAST; // @[HBMDriver.scala 92:29]
  wire [1:0] instHbm_AXI_27_RRESP; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_27_RVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_27_RREADY; // @[HBMDriver.scala 92:29]
  wire [5:0] instHbm_AXI_27_BID; // @[HBMDriver.scala 92:29]
  wire [1:0] instHbm_AXI_27_BRESP; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_27_BVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_27_BREADY; // @[HBMDriver.scala 92:29]
  wire [31:0] instHbm_AXI_27_WDATA_PARITY; // @[HBMDriver.scala 92:29]
  wire [31:0] instHbm_AXI_27_RDATA_PARITY; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_28_ACLK; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_28_ARESET_N; // @[HBMDriver.scala 92:29]
  wire [32:0] instHbm_AXI_28_ARADDR; // @[HBMDriver.scala 92:29]
  wire [1:0] instHbm_AXI_28_ARBURST; // @[HBMDriver.scala 92:29]
  wire [5:0] instHbm_AXI_28_ARID; // @[HBMDriver.scala 92:29]
  wire [3:0] instHbm_AXI_28_ARLEN; // @[HBMDriver.scala 92:29]
  wire [2:0] instHbm_AXI_28_ARSIZE; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_28_ARVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_28_ARREADY; // @[HBMDriver.scala 92:29]
  wire [32:0] instHbm_AXI_28_AWADDR; // @[HBMDriver.scala 92:29]
  wire [1:0] instHbm_AXI_28_AWBURST; // @[HBMDriver.scala 92:29]
  wire [5:0] instHbm_AXI_28_AWID; // @[HBMDriver.scala 92:29]
  wire [3:0] instHbm_AXI_28_AWLEN; // @[HBMDriver.scala 92:29]
  wire [2:0] instHbm_AXI_28_AWSIZE; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_28_AWVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_28_AWREADY; // @[HBMDriver.scala 92:29]
  wire [255:0] instHbm_AXI_28_WDATA; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_28_WLAST; // @[HBMDriver.scala 92:29]
  wire [31:0] instHbm_AXI_28_WSTRB; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_28_WVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_28_WREADY; // @[HBMDriver.scala 92:29]
  wire [255:0] instHbm_AXI_28_RDATA; // @[HBMDriver.scala 92:29]
  wire [5:0] instHbm_AXI_28_RID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_28_RLAST; // @[HBMDriver.scala 92:29]
  wire [1:0] instHbm_AXI_28_RRESP; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_28_RVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_28_RREADY; // @[HBMDriver.scala 92:29]
  wire [5:0] instHbm_AXI_28_BID; // @[HBMDriver.scala 92:29]
  wire [1:0] instHbm_AXI_28_BRESP; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_28_BVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_28_BREADY; // @[HBMDriver.scala 92:29]
  wire [31:0] instHbm_AXI_28_WDATA_PARITY; // @[HBMDriver.scala 92:29]
  wire [31:0] instHbm_AXI_28_RDATA_PARITY; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_29_ACLK; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_29_ARESET_N; // @[HBMDriver.scala 92:29]
  wire [32:0] instHbm_AXI_29_ARADDR; // @[HBMDriver.scala 92:29]
  wire [1:0] instHbm_AXI_29_ARBURST; // @[HBMDriver.scala 92:29]
  wire [5:0] instHbm_AXI_29_ARID; // @[HBMDriver.scala 92:29]
  wire [3:0] instHbm_AXI_29_ARLEN; // @[HBMDriver.scala 92:29]
  wire [2:0] instHbm_AXI_29_ARSIZE; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_29_ARVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_29_ARREADY; // @[HBMDriver.scala 92:29]
  wire [32:0] instHbm_AXI_29_AWADDR; // @[HBMDriver.scala 92:29]
  wire [1:0] instHbm_AXI_29_AWBURST; // @[HBMDriver.scala 92:29]
  wire [5:0] instHbm_AXI_29_AWID; // @[HBMDriver.scala 92:29]
  wire [3:0] instHbm_AXI_29_AWLEN; // @[HBMDriver.scala 92:29]
  wire [2:0] instHbm_AXI_29_AWSIZE; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_29_AWVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_29_AWREADY; // @[HBMDriver.scala 92:29]
  wire [255:0] instHbm_AXI_29_WDATA; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_29_WLAST; // @[HBMDriver.scala 92:29]
  wire [31:0] instHbm_AXI_29_WSTRB; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_29_WVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_29_WREADY; // @[HBMDriver.scala 92:29]
  wire [255:0] instHbm_AXI_29_RDATA; // @[HBMDriver.scala 92:29]
  wire [5:0] instHbm_AXI_29_RID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_29_RLAST; // @[HBMDriver.scala 92:29]
  wire [1:0] instHbm_AXI_29_RRESP; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_29_RVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_29_RREADY; // @[HBMDriver.scala 92:29]
  wire [5:0] instHbm_AXI_29_BID; // @[HBMDriver.scala 92:29]
  wire [1:0] instHbm_AXI_29_BRESP; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_29_BVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_29_BREADY; // @[HBMDriver.scala 92:29]
  wire [31:0] instHbm_AXI_29_WDATA_PARITY; // @[HBMDriver.scala 92:29]
  wire [31:0] instHbm_AXI_29_RDATA_PARITY; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_30_ACLK; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_30_ARESET_N; // @[HBMDriver.scala 92:29]
  wire [32:0] instHbm_AXI_30_ARADDR; // @[HBMDriver.scala 92:29]
  wire [1:0] instHbm_AXI_30_ARBURST; // @[HBMDriver.scala 92:29]
  wire [5:0] instHbm_AXI_30_ARID; // @[HBMDriver.scala 92:29]
  wire [3:0] instHbm_AXI_30_ARLEN; // @[HBMDriver.scala 92:29]
  wire [2:0] instHbm_AXI_30_ARSIZE; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_30_ARVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_30_ARREADY; // @[HBMDriver.scala 92:29]
  wire [32:0] instHbm_AXI_30_AWADDR; // @[HBMDriver.scala 92:29]
  wire [1:0] instHbm_AXI_30_AWBURST; // @[HBMDriver.scala 92:29]
  wire [5:0] instHbm_AXI_30_AWID; // @[HBMDriver.scala 92:29]
  wire [3:0] instHbm_AXI_30_AWLEN; // @[HBMDriver.scala 92:29]
  wire [2:0] instHbm_AXI_30_AWSIZE; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_30_AWVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_30_AWREADY; // @[HBMDriver.scala 92:29]
  wire [255:0] instHbm_AXI_30_WDATA; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_30_WLAST; // @[HBMDriver.scala 92:29]
  wire [31:0] instHbm_AXI_30_WSTRB; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_30_WVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_30_WREADY; // @[HBMDriver.scala 92:29]
  wire [255:0] instHbm_AXI_30_RDATA; // @[HBMDriver.scala 92:29]
  wire [5:0] instHbm_AXI_30_RID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_30_RLAST; // @[HBMDriver.scala 92:29]
  wire [1:0] instHbm_AXI_30_RRESP; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_30_RVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_30_RREADY; // @[HBMDriver.scala 92:29]
  wire [5:0] instHbm_AXI_30_BID; // @[HBMDriver.scala 92:29]
  wire [1:0] instHbm_AXI_30_BRESP; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_30_BVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_30_BREADY; // @[HBMDriver.scala 92:29]
  wire [31:0] instHbm_AXI_30_WDATA_PARITY; // @[HBMDriver.scala 92:29]
  wire [31:0] instHbm_AXI_30_RDATA_PARITY; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_31_ACLK; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_31_ARESET_N; // @[HBMDriver.scala 92:29]
  wire [32:0] instHbm_AXI_31_ARADDR; // @[HBMDriver.scala 92:29]
  wire [1:0] instHbm_AXI_31_ARBURST; // @[HBMDriver.scala 92:29]
  wire [5:0] instHbm_AXI_31_ARID; // @[HBMDriver.scala 92:29]
  wire [3:0] instHbm_AXI_31_ARLEN; // @[HBMDriver.scala 92:29]
  wire [2:0] instHbm_AXI_31_ARSIZE; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_31_ARVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_31_ARREADY; // @[HBMDriver.scala 92:29]
  wire [32:0] instHbm_AXI_31_AWADDR; // @[HBMDriver.scala 92:29]
  wire [1:0] instHbm_AXI_31_AWBURST; // @[HBMDriver.scala 92:29]
  wire [5:0] instHbm_AXI_31_AWID; // @[HBMDriver.scala 92:29]
  wire [3:0] instHbm_AXI_31_AWLEN; // @[HBMDriver.scala 92:29]
  wire [2:0] instHbm_AXI_31_AWSIZE; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_31_AWVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_31_AWREADY; // @[HBMDriver.scala 92:29]
  wire [255:0] instHbm_AXI_31_WDATA; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_31_WLAST; // @[HBMDriver.scala 92:29]
  wire [31:0] instHbm_AXI_31_WSTRB; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_31_WVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_31_WREADY; // @[HBMDriver.scala 92:29]
  wire [255:0] instHbm_AXI_31_RDATA; // @[HBMDriver.scala 92:29]
  wire [5:0] instHbm_AXI_31_RID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_31_RLAST; // @[HBMDriver.scala 92:29]
  wire [1:0] instHbm_AXI_31_RRESP; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_31_RVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_31_RREADY; // @[HBMDriver.scala 92:29]
  wire [5:0] instHbm_AXI_31_BID; // @[HBMDriver.scala 92:29]
  wire [1:0] instHbm_AXI_31_BRESP; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_31_BVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_31_BREADY; // @[HBMDriver.scala 92:29]
  wire [31:0] instHbm_AXI_31_WDATA_PARITY; // @[HBMDriver.scala 92:29]
  wire [31:0] instHbm_AXI_31_RDATA_PARITY; // @[HBMDriver.scala 92:29]
  wire [31:0] instHbm_APB_0_PWDATA; // @[HBMDriver.scala 92:29]
  wire [21:0] instHbm_APB_0_PADDR; // @[HBMDriver.scala 92:29]
  wire  instHbm_APB_0_PCLK; // @[HBMDriver.scala 92:29]
  wire  instHbm_APB_0_PENABLE; // @[HBMDriver.scala 92:29]
  wire  instHbm_APB_0_PRESET_N; // @[HBMDriver.scala 92:29]
  wire  instHbm_APB_0_PSEL; // @[HBMDriver.scala 92:29]
  wire  instHbm_APB_0_PWRITE; // @[HBMDriver.scala 92:29]
  wire [31:0] instHbm_APB_0_PRDATA; // @[HBMDriver.scala 92:29]
  wire  instHbm_APB_0_PREADY; // @[HBMDriver.scala 92:29]
  wire  instHbm_APB_0_PSLVERR; // @[HBMDriver.scala 92:29]
  wire [31:0] instHbm_APB_1_PWDATA; // @[HBMDriver.scala 92:29]
  wire [21:0] instHbm_APB_1_PADDR; // @[HBMDriver.scala 92:29]
  wire  instHbm_APB_1_PCLK; // @[HBMDriver.scala 92:29]
  wire  instHbm_APB_1_PENABLE; // @[HBMDriver.scala 92:29]
  wire  instHbm_APB_1_PRESET_N; // @[HBMDriver.scala 92:29]
  wire  instHbm_APB_1_PSEL; // @[HBMDriver.scala 92:29]
  wire  instHbm_APB_1_PWRITE; // @[HBMDriver.scala 92:29]
  wire [31:0] instHbm_APB_1_PRDATA; // @[HBMDriver.scala 92:29]
  wire  instHbm_APB_1_PREADY; // @[HBMDriver.scala 92:29]
  wire  instHbm_APB_1_PSLVERR; // @[HBMDriver.scala 92:29]
  wire  instHbm_DRAM_0_STAT_CATTRIP; // @[HBMDriver.scala 92:29]
  wire [6:0] instHbm_DRAM_0_STAT_TEMP; // @[HBMDriver.scala 92:29]
  wire  instHbm_DRAM_1_STAT_CATTRIP; // @[HBMDriver.scala 92:29]
  wire [6:0] instHbm_DRAM_1_STAT_TEMP; // @[HBMDriver.scala 92:29]
  wire  instHbm_apb_complete_0; // @[HBMDriver.scala 92:29]
  wire  instHbm_apb_complete_1; // @[HBMDriver.scala 92:29]
  reg  apb_complete_0_r; // @[Reg.scala 15:16]
  reg  apb_complete_0; // @[Reg.scala 15:16]
  reg  apb_complete_1_r; // @[Reg.scala 15:16]
  reg  apb_complete_1; // @[Reg.scala 15:16]
  reg  io_hbm_rstn_REG; // @[HBMDriver.scala 97:52]
  wire  _io_hbm_rstn_T_2 = io_hbm_rstn_REG & apb_complete_0; // @[HBMDriver.scala 98:17]
  MMCME4_ADV_Wrapper mmcmGlbl ( // @[HBMDriver.scala 48:30]
    .io_CLKIN1(mmcmGlbl_io_CLKIN1),
    .io_LOCKED(mmcmGlbl_io_LOCKED),
    .io_CLKOUT0(mmcmGlbl_io_CLKOUT0),
    .io_CLKOUT1(mmcmGlbl_io_CLKOUT1),
    .io_CLKOUT2(mmcmGlbl_io_CLKOUT2),
    .io_CLKOUT3(mmcmGlbl_io_CLKOUT3),
    .io_CLKOUT4(mmcmGlbl_io_CLKOUT4),
    .io_CLKOUT5(mmcmGlbl_io_CLKOUT5)
  );
  BUFG apb0Pclk_pad ( // @[Buf.scala 33:34]
    .O(apb0Pclk_pad_O),
    .I(apb0Pclk_pad_I)
  );
  IBUF apb0Pclk_pad_1 ( // @[Buf.scala 17:34]
    .O(apb0Pclk_pad_1_O),
    .I(apb0Pclk_pad_1_I)
  );
  BUFG apb0Pclk_pad_2 ( // @[Buf.scala 33:34]
    .O(apb0Pclk_pad_2_O),
    .I(apb0Pclk_pad_2_I)
  );
  BUFG axiAclkIn0_pad ( // @[Buf.scala 33:34]
    .O(axiAclkIn0_pad_O),
    .I(axiAclkIn0_pad_I)
  );
  BUFG hbmRefClk0_pad ( // @[Buf.scala 33:34]
    .O(hbmRefClk0_pad_O),
    .I(hbmRefClk0_pad_I)
  );
  BUFG apb1Pclk_pad ( // @[Buf.scala 33:34]
    .O(apb1Pclk_pad_O),
    .I(apb1Pclk_pad_I)
  );
  IBUF apb1Pclk_pad_1 ( // @[Buf.scala 17:34]
    .O(apb1Pclk_pad_1_O),
    .I(apb1Pclk_pad_1_I)
  );
  BUFG apb1Pclk_pad_2 ( // @[Buf.scala 33:34]
    .O(apb1Pclk_pad_2_O),
    .I(apb1Pclk_pad_2_I)
  );
  BUFG axiAclkIn1_pad ( // @[Buf.scala 33:34]
    .O(axiAclkIn1_pad_O),
    .I(axiAclkIn1_pad_I)
  );
  BUFG hbmRefClk1_pad ( // @[Buf.scala 33:34]
    .O(hbmRefClk1_pad_O),
    .I(hbmRefClk1_pad_I)
  );
  MMCME4_ADV_Wrapper_1 mmcmAxi ( // @[HBMDriver.scala 71:29]
    .io_CLKIN1(mmcmAxi_io_CLKIN1),
    .io_RST(mmcmAxi_io_RST),
    .io_LOCKED(mmcmAxi_io_LOCKED),
    .io_CLKOUT0(mmcmAxi_io_CLKOUT0)
  );
  BUFG axiAclk_pad ( // @[Buf.scala 33:34]
    .O(axiAclk_pad_O),
    .I(axiAclk_pad_I)
  );
  HBMBlackBox instHbm ( // @[HBMDriver.scala 92:29]
    .HBM_REF_CLK_0(instHbm_HBM_REF_CLK_0),
    .HBM_REF_CLK_1(instHbm_HBM_REF_CLK_1),
    .AXI_00_ACLK(instHbm_AXI_00_ACLK),
    .AXI_00_ARESET_N(instHbm_AXI_00_ARESET_N),
    .AXI_00_ARADDR(instHbm_AXI_00_ARADDR),
    .AXI_00_ARBURST(instHbm_AXI_00_ARBURST),
    .AXI_00_ARID(instHbm_AXI_00_ARID),
    .AXI_00_ARLEN(instHbm_AXI_00_ARLEN),
    .AXI_00_ARSIZE(instHbm_AXI_00_ARSIZE),
    .AXI_00_ARVALID(instHbm_AXI_00_ARVALID),
    .AXI_00_ARREADY(instHbm_AXI_00_ARREADY),
    .AXI_00_AWADDR(instHbm_AXI_00_AWADDR),
    .AXI_00_AWBURST(instHbm_AXI_00_AWBURST),
    .AXI_00_AWID(instHbm_AXI_00_AWID),
    .AXI_00_AWLEN(instHbm_AXI_00_AWLEN),
    .AXI_00_AWSIZE(instHbm_AXI_00_AWSIZE),
    .AXI_00_AWVALID(instHbm_AXI_00_AWVALID),
    .AXI_00_AWREADY(instHbm_AXI_00_AWREADY),
    .AXI_00_WDATA(instHbm_AXI_00_WDATA),
    .AXI_00_WLAST(instHbm_AXI_00_WLAST),
    .AXI_00_WSTRB(instHbm_AXI_00_WSTRB),
    .AXI_00_WVALID(instHbm_AXI_00_WVALID),
    .AXI_00_WREADY(instHbm_AXI_00_WREADY),
    .AXI_00_RDATA(instHbm_AXI_00_RDATA),
    .AXI_00_RID(instHbm_AXI_00_RID),
    .AXI_00_RLAST(instHbm_AXI_00_RLAST),
    .AXI_00_RRESP(instHbm_AXI_00_RRESP),
    .AXI_00_RVALID(instHbm_AXI_00_RVALID),
    .AXI_00_RREADY(instHbm_AXI_00_RREADY),
    .AXI_00_BID(instHbm_AXI_00_BID),
    .AXI_00_BRESP(instHbm_AXI_00_BRESP),
    .AXI_00_BVALID(instHbm_AXI_00_BVALID),
    .AXI_00_BREADY(instHbm_AXI_00_BREADY),
    .AXI_00_WDATA_PARITY(instHbm_AXI_00_WDATA_PARITY),
    .AXI_00_RDATA_PARITY(instHbm_AXI_00_RDATA_PARITY),
    .AXI_01_ACLK(instHbm_AXI_01_ACLK),
    .AXI_01_ARESET_N(instHbm_AXI_01_ARESET_N),
    .AXI_01_ARADDR(instHbm_AXI_01_ARADDR),
    .AXI_01_ARBURST(instHbm_AXI_01_ARBURST),
    .AXI_01_ARID(instHbm_AXI_01_ARID),
    .AXI_01_ARLEN(instHbm_AXI_01_ARLEN),
    .AXI_01_ARSIZE(instHbm_AXI_01_ARSIZE),
    .AXI_01_ARVALID(instHbm_AXI_01_ARVALID),
    .AXI_01_ARREADY(instHbm_AXI_01_ARREADY),
    .AXI_01_AWADDR(instHbm_AXI_01_AWADDR),
    .AXI_01_AWBURST(instHbm_AXI_01_AWBURST),
    .AXI_01_AWID(instHbm_AXI_01_AWID),
    .AXI_01_AWLEN(instHbm_AXI_01_AWLEN),
    .AXI_01_AWSIZE(instHbm_AXI_01_AWSIZE),
    .AXI_01_AWVALID(instHbm_AXI_01_AWVALID),
    .AXI_01_AWREADY(instHbm_AXI_01_AWREADY),
    .AXI_01_WDATA(instHbm_AXI_01_WDATA),
    .AXI_01_WLAST(instHbm_AXI_01_WLAST),
    .AXI_01_WSTRB(instHbm_AXI_01_WSTRB),
    .AXI_01_WVALID(instHbm_AXI_01_WVALID),
    .AXI_01_WREADY(instHbm_AXI_01_WREADY),
    .AXI_01_RDATA(instHbm_AXI_01_RDATA),
    .AXI_01_RID(instHbm_AXI_01_RID),
    .AXI_01_RLAST(instHbm_AXI_01_RLAST),
    .AXI_01_RRESP(instHbm_AXI_01_RRESP),
    .AXI_01_RVALID(instHbm_AXI_01_RVALID),
    .AXI_01_RREADY(instHbm_AXI_01_RREADY),
    .AXI_01_BID(instHbm_AXI_01_BID),
    .AXI_01_BRESP(instHbm_AXI_01_BRESP),
    .AXI_01_BVALID(instHbm_AXI_01_BVALID),
    .AXI_01_BREADY(instHbm_AXI_01_BREADY),
    .AXI_01_WDATA_PARITY(instHbm_AXI_01_WDATA_PARITY),
    .AXI_01_RDATA_PARITY(instHbm_AXI_01_RDATA_PARITY),
    .AXI_02_ACLK(instHbm_AXI_02_ACLK),
    .AXI_02_ARESET_N(instHbm_AXI_02_ARESET_N),
    .AXI_02_ARADDR(instHbm_AXI_02_ARADDR),
    .AXI_02_ARBURST(instHbm_AXI_02_ARBURST),
    .AXI_02_ARID(instHbm_AXI_02_ARID),
    .AXI_02_ARLEN(instHbm_AXI_02_ARLEN),
    .AXI_02_ARSIZE(instHbm_AXI_02_ARSIZE),
    .AXI_02_ARVALID(instHbm_AXI_02_ARVALID),
    .AXI_02_ARREADY(instHbm_AXI_02_ARREADY),
    .AXI_02_AWADDR(instHbm_AXI_02_AWADDR),
    .AXI_02_AWBURST(instHbm_AXI_02_AWBURST),
    .AXI_02_AWID(instHbm_AXI_02_AWID),
    .AXI_02_AWLEN(instHbm_AXI_02_AWLEN),
    .AXI_02_AWSIZE(instHbm_AXI_02_AWSIZE),
    .AXI_02_AWVALID(instHbm_AXI_02_AWVALID),
    .AXI_02_AWREADY(instHbm_AXI_02_AWREADY),
    .AXI_02_WDATA(instHbm_AXI_02_WDATA),
    .AXI_02_WLAST(instHbm_AXI_02_WLAST),
    .AXI_02_WSTRB(instHbm_AXI_02_WSTRB),
    .AXI_02_WVALID(instHbm_AXI_02_WVALID),
    .AXI_02_WREADY(instHbm_AXI_02_WREADY),
    .AXI_02_RDATA(instHbm_AXI_02_RDATA),
    .AXI_02_RID(instHbm_AXI_02_RID),
    .AXI_02_RLAST(instHbm_AXI_02_RLAST),
    .AXI_02_RRESP(instHbm_AXI_02_RRESP),
    .AXI_02_RVALID(instHbm_AXI_02_RVALID),
    .AXI_02_RREADY(instHbm_AXI_02_RREADY),
    .AXI_02_BID(instHbm_AXI_02_BID),
    .AXI_02_BRESP(instHbm_AXI_02_BRESP),
    .AXI_02_BVALID(instHbm_AXI_02_BVALID),
    .AXI_02_BREADY(instHbm_AXI_02_BREADY),
    .AXI_02_WDATA_PARITY(instHbm_AXI_02_WDATA_PARITY),
    .AXI_02_RDATA_PARITY(instHbm_AXI_02_RDATA_PARITY),
    .AXI_03_ACLK(instHbm_AXI_03_ACLK),
    .AXI_03_ARESET_N(instHbm_AXI_03_ARESET_N),
    .AXI_03_ARADDR(instHbm_AXI_03_ARADDR),
    .AXI_03_ARBURST(instHbm_AXI_03_ARBURST),
    .AXI_03_ARID(instHbm_AXI_03_ARID),
    .AXI_03_ARLEN(instHbm_AXI_03_ARLEN),
    .AXI_03_ARSIZE(instHbm_AXI_03_ARSIZE),
    .AXI_03_ARVALID(instHbm_AXI_03_ARVALID),
    .AXI_03_ARREADY(instHbm_AXI_03_ARREADY),
    .AXI_03_AWADDR(instHbm_AXI_03_AWADDR),
    .AXI_03_AWBURST(instHbm_AXI_03_AWBURST),
    .AXI_03_AWID(instHbm_AXI_03_AWID),
    .AXI_03_AWLEN(instHbm_AXI_03_AWLEN),
    .AXI_03_AWSIZE(instHbm_AXI_03_AWSIZE),
    .AXI_03_AWVALID(instHbm_AXI_03_AWVALID),
    .AXI_03_AWREADY(instHbm_AXI_03_AWREADY),
    .AXI_03_WDATA(instHbm_AXI_03_WDATA),
    .AXI_03_WLAST(instHbm_AXI_03_WLAST),
    .AXI_03_WSTRB(instHbm_AXI_03_WSTRB),
    .AXI_03_WVALID(instHbm_AXI_03_WVALID),
    .AXI_03_WREADY(instHbm_AXI_03_WREADY),
    .AXI_03_RDATA(instHbm_AXI_03_RDATA),
    .AXI_03_RID(instHbm_AXI_03_RID),
    .AXI_03_RLAST(instHbm_AXI_03_RLAST),
    .AXI_03_RRESP(instHbm_AXI_03_RRESP),
    .AXI_03_RVALID(instHbm_AXI_03_RVALID),
    .AXI_03_RREADY(instHbm_AXI_03_RREADY),
    .AXI_03_BID(instHbm_AXI_03_BID),
    .AXI_03_BRESP(instHbm_AXI_03_BRESP),
    .AXI_03_BVALID(instHbm_AXI_03_BVALID),
    .AXI_03_BREADY(instHbm_AXI_03_BREADY),
    .AXI_03_WDATA_PARITY(instHbm_AXI_03_WDATA_PARITY),
    .AXI_03_RDATA_PARITY(instHbm_AXI_03_RDATA_PARITY),
    .AXI_04_ACLK(instHbm_AXI_04_ACLK),
    .AXI_04_ARESET_N(instHbm_AXI_04_ARESET_N),
    .AXI_04_ARADDR(instHbm_AXI_04_ARADDR),
    .AXI_04_ARBURST(instHbm_AXI_04_ARBURST),
    .AXI_04_ARID(instHbm_AXI_04_ARID),
    .AXI_04_ARLEN(instHbm_AXI_04_ARLEN),
    .AXI_04_ARSIZE(instHbm_AXI_04_ARSIZE),
    .AXI_04_ARVALID(instHbm_AXI_04_ARVALID),
    .AXI_04_ARREADY(instHbm_AXI_04_ARREADY),
    .AXI_04_AWADDR(instHbm_AXI_04_AWADDR),
    .AXI_04_AWBURST(instHbm_AXI_04_AWBURST),
    .AXI_04_AWID(instHbm_AXI_04_AWID),
    .AXI_04_AWLEN(instHbm_AXI_04_AWLEN),
    .AXI_04_AWSIZE(instHbm_AXI_04_AWSIZE),
    .AXI_04_AWVALID(instHbm_AXI_04_AWVALID),
    .AXI_04_AWREADY(instHbm_AXI_04_AWREADY),
    .AXI_04_WDATA(instHbm_AXI_04_WDATA),
    .AXI_04_WLAST(instHbm_AXI_04_WLAST),
    .AXI_04_WSTRB(instHbm_AXI_04_WSTRB),
    .AXI_04_WVALID(instHbm_AXI_04_WVALID),
    .AXI_04_WREADY(instHbm_AXI_04_WREADY),
    .AXI_04_RDATA(instHbm_AXI_04_RDATA),
    .AXI_04_RID(instHbm_AXI_04_RID),
    .AXI_04_RLAST(instHbm_AXI_04_RLAST),
    .AXI_04_RRESP(instHbm_AXI_04_RRESP),
    .AXI_04_RVALID(instHbm_AXI_04_RVALID),
    .AXI_04_RREADY(instHbm_AXI_04_RREADY),
    .AXI_04_BID(instHbm_AXI_04_BID),
    .AXI_04_BRESP(instHbm_AXI_04_BRESP),
    .AXI_04_BVALID(instHbm_AXI_04_BVALID),
    .AXI_04_BREADY(instHbm_AXI_04_BREADY),
    .AXI_04_WDATA_PARITY(instHbm_AXI_04_WDATA_PARITY),
    .AXI_04_RDATA_PARITY(instHbm_AXI_04_RDATA_PARITY),
    .AXI_05_ACLK(instHbm_AXI_05_ACLK),
    .AXI_05_ARESET_N(instHbm_AXI_05_ARESET_N),
    .AXI_05_ARADDR(instHbm_AXI_05_ARADDR),
    .AXI_05_ARBURST(instHbm_AXI_05_ARBURST),
    .AXI_05_ARID(instHbm_AXI_05_ARID),
    .AXI_05_ARLEN(instHbm_AXI_05_ARLEN),
    .AXI_05_ARSIZE(instHbm_AXI_05_ARSIZE),
    .AXI_05_ARVALID(instHbm_AXI_05_ARVALID),
    .AXI_05_ARREADY(instHbm_AXI_05_ARREADY),
    .AXI_05_AWADDR(instHbm_AXI_05_AWADDR),
    .AXI_05_AWBURST(instHbm_AXI_05_AWBURST),
    .AXI_05_AWID(instHbm_AXI_05_AWID),
    .AXI_05_AWLEN(instHbm_AXI_05_AWLEN),
    .AXI_05_AWSIZE(instHbm_AXI_05_AWSIZE),
    .AXI_05_AWVALID(instHbm_AXI_05_AWVALID),
    .AXI_05_AWREADY(instHbm_AXI_05_AWREADY),
    .AXI_05_WDATA(instHbm_AXI_05_WDATA),
    .AXI_05_WLAST(instHbm_AXI_05_WLAST),
    .AXI_05_WSTRB(instHbm_AXI_05_WSTRB),
    .AXI_05_WVALID(instHbm_AXI_05_WVALID),
    .AXI_05_WREADY(instHbm_AXI_05_WREADY),
    .AXI_05_RDATA(instHbm_AXI_05_RDATA),
    .AXI_05_RID(instHbm_AXI_05_RID),
    .AXI_05_RLAST(instHbm_AXI_05_RLAST),
    .AXI_05_RRESP(instHbm_AXI_05_RRESP),
    .AXI_05_RVALID(instHbm_AXI_05_RVALID),
    .AXI_05_RREADY(instHbm_AXI_05_RREADY),
    .AXI_05_BID(instHbm_AXI_05_BID),
    .AXI_05_BRESP(instHbm_AXI_05_BRESP),
    .AXI_05_BVALID(instHbm_AXI_05_BVALID),
    .AXI_05_BREADY(instHbm_AXI_05_BREADY),
    .AXI_05_WDATA_PARITY(instHbm_AXI_05_WDATA_PARITY),
    .AXI_05_RDATA_PARITY(instHbm_AXI_05_RDATA_PARITY),
    .AXI_06_ACLK(instHbm_AXI_06_ACLK),
    .AXI_06_ARESET_N(instHbm_AXI_06_ARESET_N),
    .AXI_06_ARADDR(instHbm_AXI_06_ARADDR),
    .AXI_06_ARBURST(instHbm_AXI_06_ARBURST),
    .AXI_06_ARID(instHbm_AXI_06_ARID),
    .AXI_06_ARLEN(instHbm_AXI_06_ARLEN),
    .AXI_06_ARSIZE(instHbm_AXI_06_ARSIZE),
    .AXI_06_ARVALID(instHbm_AXI_06_ARVALID),
    .AXI_06_ARREADY(instHbm_AXI_06_ARREADY),
    .AXI_06_AWADDR(instHbm_AXI_06_AWADDR),
    .AXI_06_AWBURST(instHbm_AXI_06_AWBURST),
    .AXI_06_AWID(instHbm_AXI_06_AWID),
    .AXI_06_AWLEN(instHbm_AXI_06_AWLEN),
    .AXI_06_AWSIZE(instHbm_AXI_06_AWSIZE),
    .AXI_06_AWVALID(instHbm_AXI_06_AWVALID),
    .AXI_06_AWREADY(instHbm_AXI_06_AWREADY),
    .AXI_06_WDATA(instHbm_AXI_06_WDATA),
    .AXI_06_WLAST(instHbm_AXI_06_WLAST),
    .AXI_06_WSTRB(instHbm_AXI_06_WSTRB),
    .AXI_06_WVALID(instHbm_AXI_06_WVALID),
    .AXI_06_WREADY(instHbm_AXI_06_WREADY),
    .AXI_06_RDATA(instHbm_AXI_06_RDATA),
    .AXI_06_RID(instHbm_AXI_06_RID),
    .AXI_06_RLAST(instHbm_AXI_06_RLAST),
    .AXI_06_RRESP(instHbm_AXI_06_RRESP),
    .AXI_06_RVALID(instHbm_AXI_06_RVALID),
    .AXI_06_RREADY(instHbm_AXI_06_RREADY),
    .AXI_06_BID(instHbm_AXI_06_BID),
    .AXI_06_BRESP(instHbm_AXI_06_BRESP),
    .AXI_06_BVALID(instHbm_AXI_06_BVALID),
    .AXI_06_BREADY(instHbm_AXI_06_BREADY),
    .AXI_06_WDATA_PARITY(instHbm_AXI_06_WDATA_PARITY),
    .AXI_06_RDATA_PARITY(instHbm_AXI_06_RDATA_PARITY),
    .AXI_07_ACLK(instHbm_AXI_07_ACLK),
    .AXI_07_ARESET_N(instHbm_AXI_07_ARESET_N),
    .AXI_07_ARADDR(instHbm_AXI_07_ARADDR),
    .AXI_07_ARBURST(instHbm_AXI_07_ARBURST),
    .AXI_07_ARID(instHbm_AXI_07_ARID),
    .AXI_07_ARLEN(instHbm_AXI_07_ARLEN),
    .AXI_07_ARSIZE(instHbm_AXI_07_ARSIZE),
    .AXI_07_ARVALID(instHbm_AXI_07_ARVALID),
    .AXI_07_ARREADY(instHbm_AXI_07_ARREADY),
    .AXI_07_AWADDR(instHbm_AXI_07_AWADDR),
    .AXI_07_AWBURST(instHbm_AXI_07_AWBURST),
    .AXI_07_AWID(instHbm_AXI_07_AWID),
    .AXI_07_AWLEN(instHbm_AXI_07_AWLEN),
    .AXI_07_AWSIZE(instHbm_AXI_07_AWSIZE),
    .AXI_07_AWVALID(instHbm_AXI_07_AWVALID),
    .AXI_07_AWREADY(instHbm_AXI_07_AWREADY),
    .AXI_07_WDATA(instHbm_AXI_07_WDATA),
    .AXI_07_WLAST(instHbm_AXI_07_WLAST),
    .AXI_07_WSTRB(instHbm_AXI_07_WSTRB),
    .AXI_07_WVALID(instHbm_AXI_07_WVALID),
    .AXI_07_WREADY(instHbm_AXI_07_WREADY),
    .AXI_07_RDATA(instHbm_AXI_07_RDATA),
    .AXI_07_RID(instHbm_AXI_07_RID),
    .AXI_07_RLAST(instHbm_AXI_07_RLAST),
    .AXI_07_RRESP(instHbm_AXI_07_RRESP),
    .AXI_07_RVALID(instHbm_AXI_07_RVALID),
    .AXI_07_RREADY(instHbm_AXI_07_RREADY),
    .AXI_07_BID(instHbm_AXI_07_BID),
    .AXI_07_BRESP(instHbm_AXI_07_BRESP),
    .AXI_07_BVALID(instHbm_AXI_07_BVALID),
    .AXI_07_BREADY(instHbm_AXI_07_BREADY),
    .AXI_07_WDATA_PARITY(instHbm_AXI_07_WDATA_PARITY),
    .AXI_07_RDATA_PARITY(instHbm_AXI_07_RDATA_PARITY),
    .AXI_08_ACLK(instHbm_AXI_08_ACLK),
    .AXI_08_ARESET_N(instHbm_AXI_08_ARESET_N),
    .AXI_08_ARADDR(instHbm_AXI_08_ARADDR),
    .AXI_08_ARBURST(instHbm_AXI_08_ARBURST),
    .AXI_08_ARID(instHbm_AXI_08_ARID),
    .AXI_08_ARLEN(instHbm_AXI_08_ARLEN),
    .AXI_08_ARSIZE(instHbm_AXI_08_ARSIZE),
    .AXI_08_ARVALID(instHbm_AXI_08_ARVALID),
    .AXI_08_ARREADY(instHbm_AXI_08_ARREADY),
    .AXI_08_AWADDR(instHbm_AXI_08_AWADDR),
    .AXI_08_AWBURST(instHbm_AXI_08_AWBURST),
    .AXI_08_AWID(instHbm_AXI_08_AWID),
    .AXI_08_AWLEN(instHbm_AXI_08_AWLEN),
    .AXI_08_AWSIZE(instHbm_AXI_08_AWSIZE),
    .AXI_08_AWVALID(instHbm_AXI_08_AWVALID),
    .AXI_08_AWREADY(instHbm_AXI_08_AWREADY),
    .AXI_08_WDATA(instHbm_AXI_08_WDATA),
    .AXI_08_WLAST(instHbm_AXI_08_WLAST),
    .AXI_08_WSTRB(instHbm_AXI_08_WSTRB),
    .AXI_08_WVALID(instHbm_AXI_08_WVALID),
    .AXI_08_WREADY(instHbm_AXI_08_WREADY),
    .AXI_08_RDATA(instHbm_AXI_08_RDATA),
    .AXI_08_RID(instHbm_AXI_08_RID),
    .AXI_08_RLAST(instHbm_AXI_08_RLAST),
    .AXI_08_RRESP(instHbm_AXI_08_RRESP),
    .AXI_08_RVALID(instHbm_AXI_08_RVALID),
    .AXI_08_RREADY(instHbm_AXI_08_RREADY),
    .AXI_08_BID(instHbm_AXI_08_BID),
    .AXI_08_BRESP(instHbm_AXI_08_BRESP),
    .AXI_08_BVALID(instHbm_AXI_08_BVALID),
    .AXI_08_BREADY(instHbm_AXI_08_BREADY),
    .AXI_08_WDATA_PARITY(instHbm_AXI_08_WDATA_PARITY),
    .AXI_08_RDATA_PARITY(instHbm_AXI_08_RDATA_PARITY),
    .AXI_09_ACLK(instHbm_AXI_09_ACLK),
    .AXI_09_ARESET_N(instHbm_AXI_09_ARESET_N),
    .AXI_09_ARADDR(instHbm_AXI_09_ARADDR),
    .AXI_09_ARBURST(instHbm_AXI_09_ARBURST),
    .AXI_09_ARID(instHbm_AXI_09_ARID),
    .AXI_09_ARLEN(instHbm_AXI_09_ARLEN),
    .AXI_09_ARSIZE(instHbm_AXI_09_ARSIZE),
    .AXI_09_ARVALID(instHbm_AXI_09_ARVALID),
    .AXI_09_ARREADY(instHbm_AXI_09_ARREADY),
    .AXI_09_AWADDR(instHbm_AXI_09_AWADDR),
    .AXI_09_AWBURST(instHbm_AXI_09_AWBURST),
    .AXI_09_AWID(instHbm_AXI_09_AWID),
    .AXI_09_AWLEN(instHbm_AXI_09_AWLEN),
    .AXI_09_AWSIZE(instHbm_AXI_09_AWSIZE),
    .AXI_09_AWVALID(instHbm_AXI_09_AWVALID),
    .AXI_09_AWREADY(instHbm_AXI_09_AWREADY),
    .AXI_09_WDATA(instHbm_AXI_09_WDATA),
    .AXI_09_WLAST(instHbm_AXI_09_WLAST),
    .AXI_09_WSTRB(instHbm_AXI_09_WSTRB),
    .AXI_09_WVALID(instHbm_AXI_09_WVALID),
    .AXI_09_WREADY(instHbm_AXI_09_WREADY),
    .AXI_09_RDATA(instHbm_AXI_09_RDATA),
    .AXI_09_RID(instHbm_AXI_09_RID),
    .AXI_09_RLAST(instHbm_AXI_09_RLAST),
    .AXI_09_RRESP(instHbm_AXI_09_RRESP),
    .AXI_09_RVALID(instHbm_AXI_09_RVALID),
    .AXI_09_RREADY(instHbm_AXI_09_RREADY),
    .AXI_09_BID(instHbm_AXI_09_BID),
    .AXI_09_BRESP(instHbm_AXI_09_BRESP),
    .AXI_09_BVALID(instHbm_AXI_09_BVALID),
    .AXI_09_BREADY(instHbm_AXI_09_BREADY),
    .AXI_09_WDATA_PARITY(instHbm_AXI_09_WDATA_PARITY),
    .AXI_09_RDATA_PARITY(instHbm_AXI_09_RDATA_PARITY),
    .AXI_10_ACLK(instHbm_AXI_10_ACLK),
    .AXI_10_ARESET_N(instHbm_AXI_10_ARESET_N),
    .AXI_10_ARADDR(instHbm_AXI_10_ARADDR),
    .AXI_10_ARBURST(instHbm_AXI_10_ARBURST),
    .AXI_10_ARID(instHbm_AXI_10_ARID),
    .AXI_10_ARLEN(instHbm_AXI_10_ARLEN),
    .AXI_10_ARSIZE(instHbm_AXI_10_ARSIZE),
    .AXI_10_ARVALID(instHbm_AXI_10_ARVALID),
    .AXI_10_ARREADY(instHbm_AXI_10_ARREADY),
    .AXI_10_AWADDR(instHbm_AXI_10_AWADDR),
    .AXI_10_AWBURST(instHbm_AXI_10_AWBURST),
    .AXI_10_AWID(instHbm_AXI_10_AWID),
    .AXI_10_AWLEN(instHbm_AXI_10_AWLEN),
    .AXI_10_AWSIZE(instHbm_AXI_10_AWSIZE),
    .AXI_10_AWVALID(instHbm_AXI_10_AWVALID),
    .AXI_10_AWREADY(instHbm_AXI_10_AWREADY),
    .AXI_10_WDATA(instHbm_AXI_10_WDATA),
    .AXI_10_WLAST(instHbm_AXI_10_WLAST),
    .AXI_10_WSTRB(instHbm_AXI_10_WSTRB),
    .AXI_10_WVALID(instHbm_AXI_10_WVALID),
    .AXI_10_WREADY(instHbm_AXI_10_WREADY),
    .AXI_10_RDATA(instHbm_AXI_10_RDATA),
    .AXI_10_RID(instHbm_AXI_10_RID),
    .AXI_10_RLAST(instHbm_AXI_10_RLAST),
    .AXI_10_RRESP(instHbm_AXI_10_RRESP),
    .AXI_10_RVALID(instHbm_AXI_10_RVALID),
    .AXI_10_RREADY(instHbm_AXI_10_RREADY),
    .AXI_10_BID(instHbm_AXI_10_BID),
    .AXI_10_BRESP(instHbm_AXI_10_BRESP),
    .AXI_10_BVALID(instHbm_AXI_10_BVALID),
    .AXI_10_BREADY(instHbm_AXI_10_BREADY),
    .AXI_10_WDATA_PARITY(instHbm_AXI_10_WDATA_PARITY),
    .AXI_10_RDATA_PARITY(instHbm_AXI_10_RDATA_PARITY),
    .AXI_11_ACLK(instHbm_AXI_11_ACLK),
    .AXI_11_ARESET_N(instHbm_AXI_11_ARESET_N),
    .AXI_11_ARADDR(instHbm_AXI_11_ARADDR),
    .AXI_11_ARBURST(instHbm_AXI_11_ARBURST),
    .AXI_11_ARID(instHbm_AXI_11_ARID),
    .AXI_11_ARLEN(instHbm_AXI_11_ARLEN),
    .AXI_11_ARSIZE(instHbm_AXI_11_ARSIZE),
    .AXI_11_ARVALID(instHbm_AXI_11_ARVALID),
    .AXI_11_ARREADY(instHbm_AXI_11_ARREADY),
    .AXI_11_AWADDR(instHbm_AXI_11_AWADDR),
    .AXI_11_AWBURST(instHbm_AXI_11_AWBURST),
    .AXI_11_AWID(instHbm_AXI_11_AWID),
    .AXI_11_AWLEN(instHbm_AXI_11_AWLEN),
    .AXI_11_AWSIZE(instHbm_AXI_11_AWSIZE),
    .AXI_11_AWVALID(instHbm_AXI_11_AWVALID),
    .AXI_11_AWREADY(instHbm_AXI_11_AWREADY),
    .AXI_11_WDATA(instHbm_AXI_11_WDATA),
    .AXI_11_WLAST(instHbm_AXI_11_WLAST),
    .AXI_11_WSTRB(instHbm_AXI_11_WSTRB),
    .AXI_11_WVALID(instHbm_AXI_11_WVALID),
    .AXI_11_WREADY(instHbm_AXI_11_WREADY),
    .AXI_11_RDATA(instHbm_AXI_11_RDATA),
    .AXI_11_RID(instHbm_AXI_11_RID),
    .AXI_11_RLAST(instHbm_AXI_11_RLAST),
    .AXI_11_RRESP(instHbm_AXI_11_RRESP),
    .AXI_11_RVALID(instHbm_AXI_11_RVALID),
    .AXI_11_RREADY(instHbm_AXI_11_RREADY),
    .AXI_11_BID(instHbm_AXI_11_BID),
    .AXI_11_BRESP(instHbm_AXI_11_BRESP),
    .AXI_11_BVALID(instHbm_AXI_11_BVALID),
    .AXI_11_BREADY(instHbm_AXI_11_BREADY),
    .AXI_11_WDATA_PARITY(instHbm_AXI_11_WDATA_PARITY),
    .AXI_11_RDATA_PARITY(instHbm_AXI_11_RDATA_PARITY),
    .AXI_12_ACLK(instHbm_AXI_12_ACLK),
    .AXI_12_ARESET_N(instHbm_AXI_12_ARESET_N),
    .AXI_12_ARADDR(instHbm_AXI_12_ARADDR),
    .AXI_12_ARBURST(instHbm_AXI_12_ARBURST),
    .AXI_12_ARID(instHbm_AXI_12_ARID),
    .AXI_12_ARLEN(instHbm_AXI_12_ARLEN),
    .AXI_12_ARSIZE(instHbm_AXI_12_ARSIZE),
    .AXI_12_ARVALID(instHbm_AXI_12_ARVALID),
    .AXI_12_ARREADY(instHbm_AXI_12_ARREADY),
    .AXI_12_AWADDR(instHbm_AXI_12_AWADDR),
    .AXI_12_AWBURST(instHbm_AXI_12_AWBURST),
    .AXI_12_AWID(instHbm_AXI_12_AWID),
    .AXI_12_AWLEN(instHbm_AXI_12_AWLEN),
    .AXI_12_AWSIZE(instHbm_AXI_12_AWSIZE),
    .AXI_12_AWVALID(instHbm_AXI_12_AWVALID),
    .AXI_12_AWREADY(instHbm_AXI_12_AWREADY),
    .AXI_12_WDATA(instHbm_AXI_12_WDATA),
    .AXI_12_WLAST(instHbm_AXI_12_WLAST),
    .AXI_12_WSTRB(instHbm_AXI_12_WSTRB),
    .AXI_12_WVALID(instHbm_AXI_12_WVALID),
    .AXI_12_WREADY(instHbm_AXI_12_WREADY),
    .AXI_12_RDATA(instHbm_AXI_12_RDATA),
    .AXI_12_RID(instHbm_AXI_12_RID),
    .AXI_12_RLAST(instHbm_AXI_12_RLAST),
    .AXI_12_RRESP(instHbm_AXI_12_RRESP),
    .AXI_12_RVALID(instHbm_AXI_12_RVALID),
    .AXI_12_RREADY(instHbm_AXI_12_RREADY),
    .AXI_12_BID(instHbm_AXI_12_BID),
    .AXI_12_BRESP(instHbm_AXI_12_BRESP),
    .AXI_12_BVALID(instHbm_AXI_12_BVALID),
    .AXI_12_BREADY(instHbm_AXI_12_BREADY),
    .AXI_12_WDATA_PARITY(instHbm_AXI_12_WDATA_PARITY),
    .AXI_12_RDATA_PARITY(instHbm_AXI_12_RDATA_PARITY),
    .AXI_13_ACLK(instHbm_AXI_13_ACLK),
    .AXI_13_ARESET_N(instHbm_AXI_13_ARESET_N),
    .AXI_13_ARADDR(instHbm_AXI_13_ARADDR),
    .AXI_13_ARBURST(instHbm_AXI_13_ARBURST),
    .AXI_13_ARID(instHbm_AXI_13_ARID),
    .AXI_13_ARLEN(instHbm_AXI_13_ARLEN),
    .AXI_13_ARSIZE(instHbm_AXI_13_ARSIZE),
    .AXI_13_ARVALID(instHbm_AXI_13_ARVALID),
    .AXI_13_ARREADY(instHbm_AXI_13_ARREADY),
    .AXI_13_AWADDR(instHbm_AXI_13_AWADDR),
    .AXI_13_AWBURST(instHbm_AXI_13_AWBURST),
    .AXI_13_AWID(instHbm_AXI_13_AWID),
    .AXI_13_AWLEN(instHbm_AXI_13_AWLEN),
    .AXI_13_AWSIZE(instHbm_AXI_13_AWSIZE),
    .AXI_13_AWVALID(instHbm_AXI_13_AWVALID),
    .AXI_13_AWREADY(instHbm_AXI_13_AWREADY),
    .AXI_13_WDATA(instHbm_AXI_13_WDATA),
    .AXI_13_WLAST(instHbm_AXI_13_WLAST),
    .AXI_13_WSTRB(instHbm_AXI_13_WSTRB),
    .AXI_13_WVALID(instHbm_AXI_13_WVALID),
    .AXI_13_WREADY(instHbm_AXI_13_WREADY),
    .AXI_13_RDATA(instHbm_AXI_13_RDATA),
    .AXI_13_RID(instHbm_AXI_13_RID),
    .AXI_13_RLAST(instHbm_AXI_13_RLAST),
    .AXI_13_RRESP(instHbm_AXI_13_RRESP),
    .AXI_13_RVALID(instHbm_AXI_13_RVALID),
    .AXI_13_RREADY(instHbm_AXI_13_RREADY),
    .AXI_13_BID(instHbm_AXI_13_BID),
    .AXI_13_BRESP(instHbm_AXI_13_BRESP),
    .AXI_13_BVALID(instHbm_AXI_13_BVALID),
    .AXI_13_BREADY(instHbm_AXI_13_BREADY),
    .AXI_13_WDATA_PARITY(instHbm_AXI_13_WDATA_PARITY),
    .AXI_13_RDATA_PARITY(instHbm_AXI_13_RDATA_PARITY),
    .AXI_14_ACLK(instHbm_AXI_14_ACLK),
    .AXI_14_ARESET_N(instHbm_AXI_14_ARESET_N),
    .AXI_14_ARADDR(instHbm_AXI_14_ARADDR),
    .AXI_14_ARBURST(instHbm_AXI_14_ARBURST),
    .AXI_14_ARID(instHbm_AXI_14_ARID),
    .AXI_14_ARLEN(instHbm_AXI_14_ARLEN),
    .AXI_14_ARSIZE(instHbm_AXI_14_ARSIZE),
    .AXI_14_ARVALID(instHbm_AXI_14_ARVALID),
    .AXI_14_ARREADY(instHbm_AXI_14_ARREADY),
    .AXI_14_AWADDR(instHbm_AXI_14_AWADDR),
    .AXI_14_AWBURST(instHbm_AXI_14_AWBURST),
    .AXI_14_AWID(instHbm_AXI_14_AWID),
    .AXI_14_AWLEN(instHbm_AXI_14_AWLEN),
    .AXI_14_AWSIZE(instHbm_AXI_14_AWSIZE),
    .AXI_14_AWVALID(instHbm_AXI_14_AWVALID),
    .AXI_14_AWREADY(instHbm_AXI_14_AWREADY),
    .AXI_14_WDATA(instHbm_AXI_14_WDATA),
    .AXI_14_WLAST(instHbm_AXI_14_WLAST),
    .AXI_14_WSTRB(instHbm_AXI_14_WSTRB),
    .AXI_14_WVALID(instHbm_AXI_14_WVALID),
    .AXI_14_WREADY(instHbm_AXI_14_WREADY),
    .AXI_14_RDATA(instHbm_AXI_14_RDATA),
    .AXI_14_RID(instHbm_AXI_14_RID),
    .AXI_14_RLAST(instHbm_AXI_14_RLAST),
    .AXI_14_RRESP(instHbm_AXI_14_RRESP),
    .AXI_14_RVALID(instHbm_AXI_14_RVALID),
    .AXI_14_RREADY(instHbm_AXI_14_RREADY),
    .AXI_14_BID(instHbm_AXI_14_BID),
    .AXI_14_BRESP(instHbm_AXI_14_BRESP),
    .AXI_14_BVALID(instHbm_AXI_14_BVALID),
    .AXI_14_BREADY(instHbm_AXI_14_BREADY),
    .AXI_14_WDATA_PARITY(instHbm_AXI_14_WDATA_PARITY),
    .AXI_14_RDATA_PARITY(instHbm_AXI_14_RDATA_PARITY),
    .AXI_15_ACLK(instHbm_AXI_15_ACLK),
    .AXI_15_ARESET_N(instHbm_AXI_15_ARESET_N),
    .AXI_15_ARADDR(instHbm_AXI_15_ARADDR),
    .AXI_15_ARBURST(instHbm_AXI_15_ARBURST),
    .AXI_15_ARID(instHbm_AXI_15_ARID),
    .AXI_15_ARLEN(instHbm_AXI_15_ARLEN),
    .AXI_15_ARSIZE(instHbm_AXI_15_ARSIZE),
    .AXI_15_ARVALID(instHbm_AXI_15_ARVALID),
    .AXI_15_ARREADY(instHbm_AXI_15_ARREADY),
    .AXI_15_AWADDR(instHbm_AXI_15_AWADDR),
    .AXI_15_AWBURST(instHbm_AXI_15_AWBURST),
    .AXI_15_AWID(instHbm_AXI_15_AWID),
    .AXI_15_AWLEN(instHbm_AXI_15_AWLEN),
    .AXI_15_AWSIZE(instHbm_AXI_15_AWSIZE),
    .AXI_15_AWVALID(instHbm_AXI_15_AWVALID),
    .AXI_15_AWREADY(instHbm_AXI_15_AWREADY),
    .AXI_15_WDATA(instHbm_AXI_15_WDATA),
    .AXI_15_WLAST(instHbm_AXI_15_WLAST),
    .AXI_15_WSTRB(instHbm_AXI_15_WSTRB),
    .AXI_15_WVALID(instHbm_AXI_15_WVALID),
    .AXI_15_WREADY(instHbm_AXI_15_WREADY),
    .AXI_15_RDATA(instHbm_AXI_15_RDATA),
    .AXI_15_RID(instHbm_AXI_15_RID),
    .AXI_15_RLAST(instHbm_AXI_15_RLAST),
    .AXI_15_RRESP(instHbm_AXI_15_RRESP),
    .AXI_15_RVALID(instHbm_AXI_15_RVALID),
    .AXI_15_RREADY(instHbm_AXI_15_RREADY),
    .AXI_15_BID(instHbm_AXI_15_BID),
    .AXI_15_BRESP(instHbm_AXI_15_BRESP),
    .AXI_15_BVALID(instHbm_AXI_15_BVALID),
    .AXI_15_BREADY(instHbm_AXI_15_BREADY),
    .AXI_15_WDATA_PARITY(instHbm_AXI_15_WDATA_PARITY),
    .AXI_15_RDATA_PARITY(instHbm_AXI_15_RDATA_PARITY),
    .AXI_16_ACLK(instHbm_AXI_16_ACLK),
    .AXI_16_ARESET_N(instHbm_AXI_16_ARESET_N),
    .AXI_16_ARADDR(instHbm_AXI_16_ARADDR),
    .AXI_16_ARBURST(instHbm_AXI_16_ARBURST),
    .AXI_16_ARID(instHbm_AXI_16_ARID),
    .AXI_16_ARLEN(instHbm_AXI_16_ARLEN),
    .AXI_16_ARSIZE(instHbm_AXI_16_ARSIZE),
    .AXI_16_ARVALID(instHbm_AXI_16_ARVALID),
    .AXI_16_ARREADY(instHbm_AXI_16_ARREADY),
    .AXI_16_AWADDR(instHbm_AXI_16_AWADDR),
    .AXI_16_AWBURST(instHbm_AXI_16_AWBURST),
    .AXI_16_AWID(instHbm_AXI_16_AWID),
    .AXI_16_AWLEN(instHbm_AXI_16_AWLEN),
    .AXI_16_AWSIZE(instHbm_AXI_16_AWSIZE),
    .AXI_16_AWVALID(instHbm_AXI_16_AWVALID),
    .AXI_16_AWREADY(instHbm_AXI_16_AWREADY),
    .AXI_16_WDATA(instHbm_AXI_16_WDATA),
    .AXI_16_WLAST(instHbm_AXI_16_WLAST),
    .AXI_16_WSTRB(instHbm_AXI_16_WSTRB),
    .AXI_16_WVALID(instHbm_AXI_16_WVALID),
    .AXI_16_WREADY(instHbm_AXI_16_WREADY),
    .AXI_16_RDATA(instHbm_AXI_16_RDATA),
    .AXI_16_RID(instHbm_AXI_16_RID),
    .AXI_16_RLAST(instHbm_AXI_16_RLAST),
    .AXI_16_RRESP(instHbm_AXI_16_RRESP),
    .AXI_16_RVALID(instHbm_AXI_16_RVALID),
    .AXI_16_RREADY(instHbm_AXI_16_RREADY),
    .AXI_16_BID(instHbm_AXI_16_BID),
    .AXI_16_BRESP(instHbm_AXI_16_BRESP),
    .AXI_16_BVALID(instHbm_AXI_16_BVALID),
    .AXI_16_BREADY(instHbm_AXI_16_BREADY),
    .AXI_16_WDATA_PARITY(instHbm_AXI_16_WDATA_PARITY),
    .AXI_16_RDATA_PARITY(instHbm_AXI_16_RDATA_PARITY),
    .AXI_17_ACLK(instHbm_AXI_17_ACLK),
    .AXI_17_ARESET_N(instHbm_AXI_17_ARESET_N),
    .AXI_17_ARADDR(instHbm_AXI_17_ARADDR),
    .AXI_17_ARBURST(instHbm_AXI_17_ARBURST),
    .AXI_17_ARID(instHbm_AXI_17_ARID),
    .AXI_17_ARLEN(instHbm_AXI_17_ARLEN),
    .AXI_17_ARSIZE(instHbm_AXI_17_ARSIZE),
    .AXI_17_ARVALID(instHbm_AXI_17_ARVALID),
    .AXI_17_ARREADY(instHbm_AXI_17_ARREADY),
    .AXI_17_AWADDR(instHbm_AXI_17_AWADDR),
    .AXI_17_AWBURST(instHbm_AXI_17_AWBURST),
    .AXI_17_AWID(instHbm_AXI_17_AWID),
    .AXI_17_AWLEN(instHbm_AXI_17_AWLEN),
    .AXI_17_AWSIZE(instHbm_AXI_17_AWSIZE),
    .AXI_17_AWVALID(instHbm_AXI_17_AWVALID),
    .AXI_17_AWREADY(instHbm_AXI_17_AWREADY),
    .AXI_17_WDATA(instHbm_AXI_17_WDATA),
    .AXI_17_WLAST(instHbm_AXI_17_WLAST),
    .AXI_17_WSTRB(instHbm_AXI_17_WSTRB),
    .AXI_17_WVALID(instHbm_AXI_17_WVALID),
    .AXI_17_WREADY(instHbm_AXI_17_WREADY),
    .AXI_17_RDATA(instHbm_AXI_17_RDATA),
    .AXI_17_RID(instHbm_AXI_17_RID),
    .AXI_17_RLAST(instHbm_AXI_17_RLAST),
    .AXI_17_RRESP(instHbm_AXI_17_RRESP),
    .AXI_17_RVALID(instHbm_AXI_17_RVALID),
    .AXI_17_RREADY(instHbm_AXI_17_RREADY),
    .AXI_17_BID(instHbm_AXI_17_BID),
    .AXI_17_BRESP(instHbm_AXI_17_BRESP),
    .AXI_17_BVALID(instHbm_AXI_17_BVALID),
    .AXI_17_BREADY(instHbm_AXI_17_BREADY),
    .AXI_17_WDATA_PARITY(instHbm_AXI_17_WDATA_PARITY),
    .AXI_17_RDATA_PARITY(instHbm_AXI_17_RDATA_PARITY),
    .AXI_18_ACLK(instHbm_AXI_18_ACLK),
    .AXI_18_ARESET_N(instHbm_AXI_18_ARESET_N),
    .AXI_18_ARADDR(instHbm_AXI_18_ARADDR),
    .AXI_18_ARBURST(instHbm_AXI_18_ARBURST),
    .AXI_18_ARID(instHbm_AXI_18_ARID),
    .AXI_18_ARLEN(instHbm_AXI_18_ARLEN),
    .AXI_18_ARSIZE(instHbm_AXI_18_ARSIZE),
    .AXI_18_ARVALID(instHbm_AXI_18_ARVALID),
    .AXI_18_ARREADY(instHbm_AXI_18_ARREADY),
    .AXI_18_AWADDR(instHbm_AXI_18_AWADDR),
    .AXI_18_AWBURST(instHbm_AXI_18_AWBURST),
    .AXI_18_AWID(instHbm_AXI_18_AWID),
    .AXI_18_AWLEN(instHbm_AXI_18_AWLEN),
    .AXI_18_AWSIZE(instHbm_AXI_18_AWSIZE),
    .AXI_18_AWVALID(instHbm_AXI_18_AWVALID),
    .AXI_18_AWREADY(instHbm_AXI_18_AWREADY),
    .AXI_18_WDATA(instHbm_AXI_18_WDATA),
    .AXI_18_WLAST(instHbm_AXI_18_WLAST),
    .AXI_18_WSTRB(instHbm_AXI_18_WSTRB),
    .AXI_18_WVALID(instHbm_AXI_18_WVALID),
    .AXI_18_WREADY(instHbm_AXI_18_WREADY),
    .AXI_18_RDATA(instHbm_AXI_18_RDATA),
    .AXI_18_RID(instHbm_AXI_18_RID),
    .AXI_18_RLAST(instHbm_AXI_18_RLAST),
    .AXI_18_RRESP(instHbm_AXI_18_RRESP),
    .AXI_18_RVALID(instHbm_AXI_18_RVALID),
    .AXI_18_RREADY(instHbm_AXI_18_RREADY),
    .AXI_18_BID(instHbm_AXI_18_BID),
    .AXI_18_BRESP(instHbm_AXI_18_BRESP),
    .AXI_18_BVALID(instHbm_AXI_18_BVALID),
    .AXI_18_BREADY(instHbm_AXI_18_BREADY),
    .AXI_18_WDATA_PARITY(instHbm_AXI_18_WDATA_PARITY),
    .AXI_18_RDATA_PARITY(instHbm_AXI_18_RDATA_PARITY),
    .AXI_19_ACLK(instHbm_AXI_19_ACLK),
    .AXI_19_ARESET_N(instHbm_AXI_19_ARESET_N),
    .AXI_19_ARADDR(instHbm_AXI_19_ARADDR),
    .AXI_19_ARBURST(instHbm_AXI_19_ARBURST),
    .AXI_19_ARID(instHbm_AXI_19_ARID),
    .AXI_19_ARLEN(instHbm_AXI_19_ARLEN),
    .AXI_19_ARSIZE(instHbm_AXI_19_ARSIZE),
    .AXI_19_ARVALID(instHbm_AXI_19_ARVALID),
    .AXI_19_ARREADY(instHbm_AXI_19_ARREADY),
    .AXI_19_AWADDR(instHbm_AXI_19_AWADDR),
    .AXI_19_AWBURST(instHbm_AXI_19_AWBURST),
    .AXI_19_AWID(instHbm_AXI_19_AWID),
    .AXI_19_AWLEN(instHbm_AXI_19_AWLEN),
    .AXI_19_AWSIZE(instHbm_AXI_19_AWSIZE),
    .AXI_19_AWVALID(instHbm_AXI_19_AWVALID),
    .AXI_19_AWREADY(instHbm_AXI_19_AWREADY),
    .AXI_19_WDATA(instHbm_AXI_19_WDATA),
    .AXI_19_WLAST(instHbm_AXI_19_WLAST),
    .AXI_19_WSTRB(instHbm_AXI_19_WSTRB),
    .AXI_19_WVALID(instHbm_AXI_19_WVALID),
    .AXI_19_WREADY(instHbm_AXI_19_WREADY),
    .AXI_19_RDATA(instHbm_AXI_19_RDATA),
    .AXI_19_RID(instHbm_AXI_19_RID),
    .AXI_19_RLAST(instHbm_AXI_19_RLAST),
    .AXI_19_RRESP(instHbm_AXI_19_RRESP),
    .AXI_19_RVALID(instHbm_AXI_19_RVALID),
    .AXI_19_RREADY(instHbm_AXI_19_RREADY),
    .AXI_19_BID(instHbm_AXI_19_BID),
    .AXI_19_BRESP(instHbm_AXI_19_BRESP),
    .AXI_19_BVALID(instHbm_AXI_19_BVALID),
    .AXI_19_BREADY(instHbm_AXI_19_BREADY),
    .AXI_19_WDATA_PARITY(instHbm_AXI_19_WDATA_PARITY),
    .AXI_19_RDATA_PARITY(instHbm_AXI_19_RDATA_PARITY),
    .AXI_20_ACLK(instHbm_AXI_20_ACLK),
    .AXI_20_ARESET_N(instHbm_AXI_20_ARESET_N),
    .AXI_20_ARADDR(instHbm_AXI_20_ARADDR),
    .AXI_20_ARBURST(instHbm_AXI_20_ARBURST),
    .AXI_20_ARID(instHbm_AXI_20_ARID),
    .AXI_20_ARLEN(instHbm_AXI_20_ARLEN),
    .AXI_20_ARSIZE(instHbm_AXI_20_ARSIZE),
    .AXI_20_ARVALID(instHbm_AXI_20_ARVALID),
    .AXI_20_ARREADY(instHbm_AXI_20_ARREADY),
    .AXI_20_AWADDR(instHbm_AXI_20_AWADDR),
    .AXI_20_AWBURST(instHbm_AXI_20_AWBURST),
    .AXI_20_AWID(instHbm_AXI_20_AWID),
    .AXI_20_AWLEN(instHbm_AXI_20_AWLEN),
    .AXI_20_AWSIZE(instHbm_AXI_20_AWSIZE),
    .AXI_20_AWVALID(instHbm_AXI_20_AWVALID),
    .AXI_20_AWREADY(instHbm_AXI_20_AWREADY),
    .AXI_20_WDATA(instHbm_AXI_20_WDATA),
    .AXI_20_WLAST(instHbm_AXI_20_WLAST),
    .AXI_20_WSTRB(instHbm_AXI_20_WSTRB),
    .AXI_20_WVALID(instHbm_AXI_20_WVALID),
    .AXI_20_WREADY(instHbm_AXI_20_WREADY),
    .AXI_20_RDATA(instHbm_AXI_20_RDATA),
    .AXI_20_RID(instHbm_AXI_20_RID),
    .AXI_20_RLAST(instHbm_AXI_20_RLAST),
    .AXI_20_RRESP(instHbm_AXI_20_RRESP),
    .AXI_20_RVALID(instHbm_AXI_20_RVALID),
    .AXI_20_RREADY(instHbm_AXI_20_RREADY),
    .AXI_20_BID(instHbm_AXI_20_BID),
    .AXI_20_BRESP(instHbm_AXI_20_BRESP),
    .AXI_20_BVALID(instHbm_AXI_20_BVALID),
    .AXI_20_BREADY(instHbm_AXI_20_BREADY),
    .AXI_20_WDATA_PARITY(instHbm_AXI_20_WDATA_PARITY),
    .AXI_20_RDATA_PARITY(instHbm_AXI_20_RDATA_PARITY),
    .AXI_21_ACLK(instHbm_AXI_21_ACLK),
    .AXI_21_ARESET_N(instHbm_AXI_21_ARESET_N),
    .AXI_21_ARADDR(instHbm_AXI_21_ARADDR),
    .AXI_21_ARBURST(instHbm_AXI_21_ARBURST),
    .AXI_21_ARID(instHbm_AXI_21_ARID),
    .AXI_21_ARLEN(instHbm_AXI_21_ARLEN),
    .AXI_21_ARSIZE(instHbm_AXI_21_ARSIZE),
    .AXI_21_ARVALID(instHbm_AXI_21_ARVALID),
    .AXI_21_ARREADY(instHbm_AXI_21_ARREADY),
    .AXI_21_AWADDR(instHbm_AXI_21_AWADDR),
    .AXI_21_AWBURST(instHbm_AXI_21_AWBURST),
    .AXI_21_AWID(instHbm_AXI_21_AWID),
    .AXI_21_AWLEN(instHbm_AXI_21_AWLEN),
    .AXI_21_AWSIZE(instHbm_AXI_21_AWSIZE),
    .AXI_21_AWVALID(instHbm_AXI_21_AWVALID),
    .AXI_21_AWREADY(instHbm_AXI_21_AWREADY),
    .AXI_21_WDATA(instHbm_AXI_21_WDATA),
    .AXI_21_WLAST(instHbm_AXI_21_WLAST),
    .AXI_21_WSTRB(instHbm_AXI_21_WSTRB),
    .AXI_21_WVALID(instHbm_AXI_21_WVALID),
    .AXI_21_WREADY(instHbm_AXI_21_WREADY),
    .AXI_21_RDATA(instHbm_AXI_21_RDATA),
    .AXI_21_RID(instHbm_AXI_21_RID),
    .AXI_21_RLAST(instHbm_AXI_21_RLAST),
    .AXI_21_RRESP(instHbm_AXI_21_RRESP),
    .AXI_21_RVALID(instHbm_AXI_21_RVALID),
    .AXI_21_RREADY(instHbm_AXI_21_RREADY),
    .AXI_21_BID(instHbm_AXI_21_BID),
    .AXI_21_BRESP(instHbm_AXI_21_BRESP),
    .AXI_21_BVALID(instHbm_AXI_21_BVALID),
    .AXI_21_BREADY(instHbm_AXI_21_BREADY),
    .AXI_21_WDATA_PARITY(instHbm_AXI_21_WDATA_PARITY),
    .AXI_21_RDATA_PARITY(instHbm_AXI_21_RDATA_PARITY),
    .AXI_22_ACLK(instHbm_AXI_22_ACLK),
    .AXI_22_ARESET_N(instHbm_AXI_22_ARESET_N),
    .AXI_22_ARADDR(instHbm_AXI_22_ARADDR),
    .AXI_22_ARBURST(instHbm_AXI_22_ARBURST),
    .AXI_22_ARID(instHbm_AXI_22_ARID),
    .AXI_22_ARLEN(instHbm_AXI_22_ARLEN),
    .AXI_22_ARSIZE(instHbm_AXI_22_ARSIZE),
    .AXI_22_ARVALID(instHbm_AXI_22_ARVALID),
    .AXI_22_ARREADY(instHbm_AXI_22_ARREADY),
    .AXI_22_AWADDR(instHbm_AXI_22_AWADDR),
    .AXI_22_AWBURST(instHbm_AXI_22_AWBURST),
    .AXI_22_AWID(instHbm_AXI_22_AWID),
    .AXI_22_AWLEN(instHbm_AXI_22_AWLEN),
    .AXI_22_AWSIZE(instHbm_AXI_22_AWSIZE),
    .AXI_22_AWVALID(instHbm_AXI_22_AWVALID),
    .AXI_22_AWREADY(instHbm_AXI_22_AWREADY),
    .AXI_22_WDATA(instHbm_AXI_22_WDATA),
    .AXI_22_WLAST(instHbm_AXI_22_WLAST),
    .AXI_22_WSTRB(instHbm_AXI_22_WSTRB),
    .AXI_22_WVALID(instHbm_AXI_22_WVALID),
    .AXI_22_WREADY(instHbm_AXI_22_WREADY),
    .AXI_22_RDATA(instHbm_AXI_22_RDATA),
    .AXI_22_RID(instHbm_AXI_22_RID),
    .AXI_22_RLAST(instHbm_AXI_22_RLAST),
    .AXI_22_RRESP(instHbm_AXI_22_RRESP),
    .AXI_22_RVALID(instHbm_AXI_22_RVALID),
    .AXI_22_RREADY(instHbm_AXI_22_RREADY),
    .AXI_22_BID(instHbm_AXI_22_BID),
    .AXI_22_BRESP(instHbm_AXI_22_BRESP),
    .AXI_22_BVALID(instHbm_AXI_22_BVALID),
    .AXI_22_BREADY(instHbm_AXI_22_BREADY),
    .AXI_22_WDATA_PARITY(instHbm_AXI_22_WDATA_PARITY),
    .AXI_22_RDATA_PARITY(instHbm_AXI_22_RDATA_PARITY),
    .AXI_23_ACLK(instHbm_AXI_23_ACLK),
    .AXI_23_ARESET_N(instHbm_AXI_23_ARESET_N),
    .AXI_23_ARADDR(instHbm_AXI_23_ARADDR),
    .AXI_23_ARBURST(instHbm_AXI_23_ARBURST),
    .AXI_23_ARID(instHbm_AXI_23_ARID),
    .AXI_23_ARLEN(instHbm_AXI_23_ARLEN),
    .AXI_23_ARSIZE(instHbm_AXI_23_ARSIZE),
    .AXI_23_ARVALID(instHbm_AXI_23_ARVALID),
    .AXI_23_ARREADY(instHbm_AXI_23_ARREADY),
    .AXI_23_AWADDR(instHbm_AXI_23_AWADDR),
    .AXI_23_AWBURST(instHbm_AXI_23_AWBURST),
    .AXI_23_AWID(instHbm_AXI_23_AWID),
    .AXI_23_AWLEN(instHbm_AXI_23_AWLEN),
    .AXI_23_AWSIZE(instHbm_AXI_23_AWSIZE),
    .AXI_23_AWVALID(instHbm_AXI_23_AWVALID),
    .AXI_23_AWREADY(instHbm_AXI_23_AWREADY),
    .AXI_23_WDATA(instHbm_AXI_23_WDATA),
    .AXI_23_WLAST(instHbm_AXI_23_WLAST),
    .AXI_23_WSTRB(instHbm_AXI_23_WSTRB),
    .AXI_23_WVALID(instHbm_AXI_23_WVALID),
    .AXI_23_WREADY(instHbm_AXI_23_WREADY),
    .AXI_23_RDATA(instHbm_AXI_23_RDATA),
    .AXI_23_RID(instHbm_AXI_23_RID),
    .AXI_23_RLAST(instHbm_AXI_23_RLAST),
    .AXI_23_RRESP(instHbm_AXI_23_RRESP),
    .AXI_23_RVALID(instHbm_AXI_23_RVALID),
    .AXI_23_RREADY(instHbm_AXI_23_RREADY),
    .AXI_23_BID(instHbm_AXI_23_BID),
    .AXI_23_BRESP(instHbm_AXI_23_BRESP),
    .AXI_23_BVALID(instHbm_AXI_23_BVALID),
    .AXI_23_BREADY(instHbm_AXI_23_BREADY),
    .AXI_23_WDATA_PARITY(instHbm_AXI_23_WDATA_PARITY),
    .AXI_23_RDATA_PARITY(instHbm_AXI_23_RDATA_PARITY),
    .AXI_24_ACLK(instHbm_AXI_24_ACLK),
    .AXI_24_ARESET_N(instHbm_AXI_24_ARESET_N),
    .AXI_24_ARADDR(instHbm_AXI_24_ARADDR),
    .AXI_24_ARBURST(instHbm_AXI_24_ARBURST),
    .AXI_24_ARID(instHbm_AXI_24_ARID),
    .AXI_24_ARLEN(instHbm_AXI_24_ARLEN),
    .AXI_24_ARSIZE(instHbm_AXI_24_ARSIZE),
    .AXI_24_ARVALID(instHbm_AXI_24_ARVALID),
    .AXI_24_ARREADY(instHbm_AXI_24_ARREADY),
    .AXI_24_AWADDR(instHbm_AXI_24_AWADDR),
    .AXI_24_AWBURST(instHbm_AXI_24_AWBURST),
    .AXI_24_AWID(instHbm_AXI_24_AWID),
    .AXI_24_AWLEN(instHbm_AXI_24_AWLEN),
    .AXI_24_AWSIZE(instHbm_AXI_24_AWSIZE),
    .AXI_24_AWVALID(instHbm_AXI_24_AWVALID),
    .AXI_24_AWREADY(instHbm_AXI_24_AWREADY),
    .AXI_24_WDATA(instHbm_AXI_24_WDATA),
    .AXI_24_WLAST(instHbm_AXI_24_WLAST),
    .AXI_24_WSTRB(instHbm_AXI_24_WSTRB),
    .AXI_24_WVALID(instHbm_AXI_24_WVALID),
    .AXI_24_WREADY(instHbm_AXI_24_WREADY),
    .AXI_24_RDATA(instHbm_AXI_24_RDATA),
    .AXI_24_RID(instHbm_AXI_24_RID),
    .AXI_24_RLAST(instHbm_AXI_24_RLAST),
    .AXI_24_RRESP(instHbm_AXI_24_RRESP),
    .AXI_24_RVALID(instHbm_AXI_24_RVALID),
    .AXI_24_RREADY(instHbm_AXI_24_RREADY),
    .AXI_24_BID(instHbm_AXI_24_BID),
    .AXI_24_BRESP(instHbm_AXI_24_BRESP),
    .AXI_24_BVALID(instHbm_AXI_24_BVALID),
    .AXI_24_BREADY(instHbm_AXI_24_BREADY),
    .AXI_24_WDATA_PARITY(instHbm_AXI_24_WDATA_PARITY),
    .AXI_24_RDATA_PARITY(instHbm_AXI_24_RDATA_PARITY),
    .AXI_25_ACLK(instHbm_AXI_25_ACLK),
    .AXI_25_ARESET_N(instHbm_AXI_25_ARESET_N),
    .AXI_25_ARADDR(instHbm_AXI_25_ARADDR),
    .AXI_25_ARBURST(instHbm_AXI_25_ARBURST),
    .AXI_25_ARID(instHbm_AXI_25_ARID),
    .AXI_25_ARLEN(instHbm_AXI_25_ARLEN),
    .AXI_25_ARSIZE(instHbm_AXI_25_ARSIZE),
    .AXI_25_ARVALID(instHbm_AXI_25_ARVALID),
    .AXI_25_ARREADY(instHbm_AXI_25_ARREADY),
    .AXI_25_AWADDR(instHbm_AXI_25_AWADDR),
    .AXI_25_AWBURST(instHbm_AXI_25_AWBURST),
    .AXI_25_AWID(instHbm_AXI_25_AWID),
    .AXI_25_AWLEN(instHbm_AXI_25_AWLEN),
    .AXI_25_AWSIZE(instHbm_AXI_25_AWSIZE),
    .AXI_25_AWVALID(instHbm_AXI_25_AWVALID),
    .AXI_25_AWREADY(instHbm_AXI_25_AWREADY),
    .AXI_25_WDATA(instHbm_AXI_25_WDATA),
    .AXI_25_WLAST(instHbm_AXI_25_WLAST),
    .AXI_25_WSTRB(instHbm_AXI_25_WSTRB),
    .AXI_25_WVALID(instHbm_AXI_25_WVALID),
    .AXI_25_WREADY(instHbm_AXI_25_WREADY),
    .AXI_25_RDATA(instHbm_AXI_25_RDATA),
    .AXI_25_RID(instHbm_AXI_25_RID),
    .AXI_25_RLAST(instHbm_AXI_25_RLAST),
    .AXI_25_RRESP(instHbm_AXI_25_RRESP),
    .AXI_25_RVALID(instHbm_AXI_25_RVALID),
    .AXI_25_RREADY(instHbm_AXI_25_RREADY),
    .AXI_25_BID(instHbm_AXI_25_BID),
    .AXI_25_BRESP(instHbm_AXI_25_BRESP),
    .AXI_25_BVALID(instHbm_AXI_25_BVALID),
    .AXI_25_BREADY(instHbm_AXI_25_BREADY),
    .AXI_25_WDATA_PARITY(instHbm_AXI_25_WDATA_PARITY),
    .AXI_25_RDATA_PARITY(instHbm_AXI_25_RDATA_PARITY),
    .AXI_26_ACLK(instHbm_AXI_26_ACLK),
    .AXI_26_ARESET_N(instHbm_AXI_26_ARESET_N),
    .AXI_26_ARADDR(instHbm_AXI_26_ARADDR),
    .AXI_26_ARBURST(instHbm_AXI_26_ARBURST),
    .AXI_26_ARID(instHbm_AXI_26_ARID),
    .AXI_26_ARLEN(instHbm_AXI_26_ARLEN),
    .AXI_26_ARSIZE(instHbm_AXI_26_ARSIZE),
    .AXI_26_ARVALID(instHbm_AXI_26_ARVALID),
    .AXI_26_ARREADY(instHbm_AXI_26_ARREADY),
    .AXI_26_AWADDR(instHbm_AXI_26_AWADDR),
    .AXI_26_AWBURST(instHbm_AXI_26_AWBURST),
    .AXI_26_AWID(instHbm_AXI_26_AWID),
    .AXI_26_AWLEN(instHbm_AXI_26_AWLEN),
    .AXI_26_AWSIZE(instHbm_AXI_26_AWSIZE),
    .AXI_26_AWVALID(instHbm_AXI_26_AWVALID),
    .AXI_26_AWREADY(instHbm_AXI_26_AWREADY),
    .AXI_26_WDATA(instHbm_AXI_26_WDATA),
    .AXI_26_WLAST(instHbm_AXI_26_WLAST),
    .AXI_26_WSTRB(instHbm_AXI_26_WSTRB),
    .AXI_26_WVALID(instHbm_AXI_26_WVALID),
    .AXI_26_WREADY(instHbm_AXI_26_WREADY),
    .AXI_26_RDATA(instHbm_AXI_26_RDATA),
    .AXI_26_RID(instHbm_AXI_26_RID),
    .AXI_26_RLAST(instHbm_AXI_26_RLAST),
    .AXI_26_RRESP(instHbm_AXI_26_RRESP),
    .AXI_26_RVALID(instHbm_AXI_26_RVALID),
    .AXI_26_RREADY(instHbm_AXI_26_RREADY),
    .AXI_26_BID(instHbm_AXI_26_BID),
    .AXI_26_BRESP(instHbm_AXI_26_BRESP),
    .AXI_26_BVALID(instHbm_AXI_26_BVALID),
    .AXI_26_BREADY(instHbm_AXI_26_BREADY),
    .AXI_26_WDATA_PARITY(instHbm_AXI_26_WDATA_PARITY),
    .AXI_26_RDATA_PARITY(instHbm_AXI_26_RDATA_PARITY),
    .AXI_27_ACLK(instHbm_AXI_27_ACLK),
    .AXI_27_ARESET_N(instHbm_AXI_27_ARESET_N),
    .AXI_27_ARADDR(instHbm_AXI_27_ARADDR),
    .AXI_27_ARBURST(instHbm_AXI_27_ARBURST),
    .AXI_27_ARID(instHbm_AXI_27_ARID),
    .AXI_27_ARLEN(instHbm_AXI_27_ARLEN),
    .AXI_27_ARSIZE(instHbm_AXI_27_ARSIZE),
    .AXI_27_ARVALID(instHbm_AXI_27_ARVALID),
    .AXI_27_ARREADY(instHbm_AXI_27_ARREADY),
    .AXI_27_AWADDR(instHbm_AXI_27_AWADDR),
    .AXI_27_AWBURST(instHbm_AXI_27_AWBURST),
    .AXI_27_AWID(instHbm_AXI_27_AWID),
    .AXI_27_AWLEN(instHbm_AXI_27_AWLEN),
    .AXI_27_AWSIZE(instHbm_AXI_27_AWSIZE),
    .AXI_27_AWVALID(instHbm_AXI_27_AWVALID),
    .AXI_27_AWREADY(instHbm_AXI_27_AWREADY),
    .AXI_27_WDATA(instHbm_AXI_27_WDATA),
    .AXI_27_WLAST(instHbm_AXI_27_WLAST),
    .AXI_27_WSTRB(instHbm_AXI_27_WSTRB),
    .AXI_27_WVALID(instHbm_AXI_27_WVALID),
    .AXI_27_WREADY(instHbm_AXI_27_WREADY),
    .AXI_27_RDATA(instHbm_AXI_27_RDATA),
    .AXI_27_RID(instHbm_AXI_27_RID),
    .AXI_27_RLAST(instHbm_AXI_27_RLAST),
    .AXI_27_RRESP(instHbm_AXI_27_RRESP),
    .AXI_27_RVALID(instHbm_AXI_27_RVALID),
    .AXI_27_RREADY(instHbm_AXI_27_RREADY),
    .AXI_27_BID(instHbm_AXI_27_BID),
    .AXI_27_BRESP(instHbm_AXI_27_BRESP),
    .AXI_27_BVALID(instHbm_AXI_27_BVALID),
    .AXI_27_BREADY(instHbm_AXI_27_BREADY),
    .AXI_27_WDATA_PARITY(instHbm_AXI_27_WDATA_PARITY),
    .AXI_27_RDATA_PARITY(instHbm_AXI_27_RDATA_PARITY),
    .AXI_28_ACLK(instHbm_AXI_28_ACLK),
    .AXI_28_ARESET_N(instHbm_AXI_28_ARESET_N),
    .AXI_28_ARADDR(instHbm_AXI_28_ARADDR),
    .AXI_28_ARBURST(instHbm_AXI_28_ARBURST),
    .AXI_28_ARID(instHbm_AXI_28_ARID),
    .AXI_28_ARLEN(instHbm_AXI_28_ARLEN),
    .AXI_28_ARSIZE(instHbm_AXI_28_ARSIZE),
    .AXI_28_ARVALID(instHbm_AXI_28_ARVALID),
    .AXI_28_ARREADY(instHbm_AXI_28_ARREADY),
    .AXI_28_AWADDR(instHbm_AXI_28_AWADDR),
    .AXI_28_AWBURST(instHbm_AXI_28_AWBURST),
    .AXI_28_AWID(instHbm_AXI_28_AWID),
    .AXI_28_AWLEN(instHbm_AXI_28_AWLEN),
    .AXI_28_AWSIZE(instHbm_AXI_28_AWSIZE),
    .AXI_28_AWVALID(instHbm_AXI_28_AWVALID),
    .AXI_28_AWREADY(instHbm_AXI_28_AWREADY),
    .AXI_28_WDATA(instHbm_AXI_28_WDATA),
    .AXI_28_WLAST(instHbm_AXI_28_WLAST),
    .AXI_28_WSTRB(instHbm_AXI_28_WSTRB),
    .AXI_28_WVALID(instHbm_AXI_28_WVALID),
    .AXI_28_WREADY(instHbm_AXI_28_WREADY),
    .AXI_28_RDATA(instHbm_AXI_28_RDATA),
    .AXI_28_RID(instHbm_AXI_28_RID),
    .AXI_28_RLAST(instHbm_AXI_28_RLAST),
    .AXI_28_RRESP(instHbm_AXI_28_RRESP),
    .AXI_28_RVALID(instHbm_AXI_28_RVALID),
    .AXI_28_RREADY(instHbm_AXI_28_RREADY),
    .AXI_28_BID(instHbm_AXI_28_BID),
    .AXI_28_BRESP(instHbm_AXI_28_BRESP),
    .AXI_28_BVALID(instHbm_AXI_28_BVALID),
    .AXI_28_BREADY(instHbm_AXI_28_BREADY),
    .AXI_28_WDATA_PARITY(instHbm_AXI_28_WDATA_PARITY),
    .AXI_28_RDATA_PARITY(instHbm_AXI_28_RDATA_PARITY),
    .AXI_29_ACLK(instHbm_AXI_29_ACLK),
    .AXI_29_ARESET_N(instHbm_AXI_29_ARESET_N),
    .AXI_29_ARADDR(instHbm_AXI_29_ARADDR),
    .AXI_29_ARBURST(instHbm_AXI_29_ARBURST),
    .AXI_29_ARID(instHbm_AXI_29_ARID),
    .AXI_29_ARLEN(instHbm_AXI_29_ARLEN),
    .AXI_29_ARSIZE(instHbm_AXI_29_ARSIZE),
    .AXI_29_ARVALID(instHbm_AXI_29_ARVALID),
    .AXI_29_ARREADY(instHbm_AXI_29_ARREADY),
    .AXI_29_AWADDR(instHbm_AXI_29_AWADDR),
    .AXI_29_AWBURST(instHbm_AXI_29_AWBURST),
    .AXI_29_AWID(instHbm_AXI_29_AWID),
    .AXI_29_AWLEN(instHbm_AXI_29_AWLEN),
    .AXI_29_AWSIZE(instHbm_AXI_29_AWSIZE),
    .AXI_29_AWVALID(instHbm_AXI_29_AWVALID),
    .AXI_29_AWREADY(instHbm_AXI_29_AWREADY),
    .AXI_29_WDATA(instHbm_AXI_29_WDATA),
    .AXI_29_WLAST(instHbm_AXI_29_WLAST),
    .AXI_29_WSTRB(instHbm_AXI_29_WSTRB),
    .AXI_29_WVALID(instHbm_AXI_29_WVALID),
    .AXI_29_WREADY(instHbm_AXI_29_WREADY),
    .AXI_29_RDATA(instHbm_AXI_29_RDATA),
    .AXI_29_RID(instHbm_AXI_29_RID),
    .AXI_29_RLAST(instHbm_AXI_29_RLAST),
    .AXI_29_RRESP(instHbm_AXI_29_RRESP),
    .AXI_29_RVALID(instHbm_AXI_29_RVALID),
    .AXI_29_RREADY(instHbm_AXI_29_RREADY),
    .AXI_29_BID(instHbm_AXI_29_BID),
    .AXI_29_BRESP(instHbm_AXI_29_BRESP),
    .AXI_29_BVALID(instHbm_AXI_29_BVALID),
    .AXI_29_BREADY(instHbm_AXI_29_BREADY),
    .AXI_29_WDATA_PARITY(instHbm_AXI_29_WDATA_PARITY),
    .AXI_29_RDATA_PARITY(instHbm_AXI_29_RDATA_PARITY),
    .AXI_30_ACLK(instHbm_AXI_30_ACLK),
    .AXI_30_ARESET_N(instHbm_AXI_30_ARESET_N),
    .AXI_30_ARADDR(instHbm_AXI_30_ARADDR),
    .AXI_30_ARBURST(instHbm_AXI_30_ARBURST),
    .AXI_30_ARID(instHbm_AXI_30_ARID),
    .AXI_30_ARLEN(instHbm_AXI_30_ARLEN),
    .AXI_30_ARSIZE(instHbm_AXI_30_ARSIZE),
    .AXI_30_ARVALID(instHbm_AXI_30_ARVALID),
    .AXI_30_ARREADY(instHbm_AXI_30_ARREADY),
    .AXI_30_AWADDR(instHbm_AXI_30_AWADDR),
    .AXI_30_AWBURST(instHbm_AXI_30_AWBURST),
    .AXI_30_AWID(instHbm_AXI_30_AWID),
    .AXI_30_AWLEN(instHbm_AXI_30_AWLEN),
    .AXI_30_AWSIZE(instHbm_AXI_30_AWSIZE),
    .AXI_30_AWVALID(instHbm_AXI_30_AWVALID),
    .AXI_30_AWREADY(instHbm_AXI_30_AWREADY),
    .AXI_30_WDATA(instHbm_AXI_30_WDATA),
    .AXI_30_WLAST(instHbm_AXI_30_WLAST),
    .AXI_30_WSTRB(instHbm_AXI_30_WSTRB),
    .AXI_30_WVALID(instHbm_AXI_30_WVALID),
    .AXI_30_WREADY(instHbm_AXI_30_WREADY),
    .AXI_30_RDATA(instHbm_AXI_30_RDATA),
    .AXI_30_RID(instHbm_AXI_30_RID),
    .AXI_30_RLAST(instHbm_AXI_30_RLAST),
    .AXI_30_RRESP(instHbm_AXI_30_RRESP),
    .AXI_30_RVALID(instHbm_AXI_30_RVALID),
    .AXI_30_RREADY(instHbm_AXI_30_RREADY),
    .AXI_30_BID(instHbm_AXI_30_BID),
    .AXI_30_BRESP(instHbm_AXI_30_BRESP),
    .AXI_30_BVALID(instHbm_AXI_30_BVALID),
    .AXI_30_BREADY(instHbm_AXI_30_BREADY),
    .AXI_30_WDATA_PARITY(instHbm_AXI_30_WDATA_PARITY),
    .AXI_30_RDATA_PARITY(instHbm_AXI_30_RDATA_PARITY),
    .AXI_31_ACLK(instHbm_AXI_31_ACLK),
    .AXI_31_ARESET_N(instHbm_AXI_31_ARESET_N),
    .AXI_31_ARADDR(instHbm_AXI_31_ARADDR),
    .AXI_31_ARBURST(instHbm_AXI_31_ARBURST),
    .AXI_31_ARID(instHbm_AXI_31_ARID),
    .AXI_31_ARLEN(instHbm_AXI_31_ARLEN),
    .AXI_31_ARSIZE(instHbm_AXI_31_ARSIZE),
    .AXI_31_ARVALID(instHbm_AXI_31_ARVALID),
    .AXI_31_ARREADY(instHbm_AXI_31_ARREADY),
    .AXI_31_AWADDR(instHbm_AXI_31_AWADDR),
    .AXI_31_AWBURST(instHbm_AXI_31_AWBURST),
    .AXI_31_AWID(instHbm_AXI_31_AWID),
    .AXI_31_AWLEN(instHbm_AXI_31_AWLEN),
    .AXI_31_AWSIZE(instHbm_AXI_31_AWSIZE),
    .AXI_31_AWVALID(instHbm_AXI_31_AWVALID),
    .AXI_31_AWREADY(instHbm_AXI_31_AWREADY),
    .AXI_31_WDATA(instHbm_AXI_31_WDATA),
    .AXI_31_WLAST(instHbm_AXI_31_WLAST),
    .AXI_31_WSTRB(instHbm_AXI_31_WSTRB),
    .AXI_31_WVALID(instHbm_AXI_31_WVALID),
    .AXI_31_WREADY(instHbm_AXI_31_WREADY),
    .AXI_31_RDATA(instHbm_AXI_31_RDATA),
    .AXI_31_RID(instHbm_AXI_31_RID),
    .AXI_31_RLAST(instHbm_AXI_31_RLAST),
    .AXI_31_RRESP(instHbm_AXI_31_RRESP),
    .AXI_31_RVALID(instHbm_AXI_31_RVALID),
    .AXI_31_RREADY(instHbm_AXI_31_RREADY),
    .AXI_31_BID(instHbm_AXI_31_BID),
    .AXI_31_BRESP(instHbm_AXI_31_BRESP),
    .AXI_31_BVALID(instHbm_AXI_31_BVALID),
    .AXI_31_BREADY(instHbm_AXI_31_BREADY),
    .AXI_31_WDATA_PARITY(instHbm_AXI_31_WDATA_PARITY),
    .AXI_31_RDATA_PARITY(instHbm_AXI_31_RDATA_PARITY),
    .APB_0_PWDATA(instHbm_APB_0_PWDATA),
    .APB_0_PADDR(instHbm_APB_0_PADDR),
    .APB_0_PCLK(instHbm_APB_0_PCLK),
    .APB_0_PENABLE(instHbm_APB_0_PENABLE),
    .APB_0_PRESET_N(instHbm_APB_0_PRESET_N),
    .APB_0_PSEL(instHbm_APB_0_PSEL),
    .APB_0_PWRITE(instHbm_APB_0_PWRITE),
    .APB_0_PRDATA(instHbm_APB_0_PRDATA),
    .APB_0_PREADY(instHbm_APB_0_PREADY),
    .APB_0_PSLVERR(instHbm_APB_0_PSLVERR),
    .APB_1_PWDATA(instHbm_APB_1_PWDATA),
    .APB_1_PADDR(instHbm_APB_1_PADDR),
    .APB_1_PCLK(instHbm_APB_1_PCLK),
    .APB_1_PENABLE(instHbm_APB_1_PENABLE),
    .APB_1_PRESET_N(instHbm_APB_1_PRESET_N),
    .APB_1_PSEL(instHbm_APB_1_PSEL),
    .APB_1_PWRITE(instHbm_APB_1_PWRITE),
    .APB_1_PRDATA(instHbm_APB_1_PRDATA),
    .APB_1_PREADY(instHbm_APB_1_PREADY),
    .APB_1_PSLVERR(instHbm_APB_1_PSLVERR),
    .DRAM_0_STAT_CATTRIP(instHbm_DRAM_0_STAT_CATTRIP),
    .DRAM_0_STAT_TEMP(instHbm_DRAM_0_STAT_TEMP),
    .DRAM_1_STAT_CATTRIP(instHbm_DRAM_1_STAT_CATTRIP),
    .DRAM_1_STAT_TEMP(instHbm_DRAM_1_STAT_TEMP),
    .apb_complete_0(instHbm_apb_complete_0),
    .apb_complete_1(instHbm_apb_complete_1)
  );
  assign io_hbm_clk = axiAclk_pad_O; // @[HBMDriver.scala 90:25]
  assign io_hbm_rstn = _io_hbm_rstn_T_2 & apb_complete_1; // @[HBMDriver.scala 99:17]
  assign mmcmGlbl_io_CLKIN1 = clock; // @[HBMDriver.scala 60:33]
  assign apb0Pclk_pad_I = mmcmGlbl_io_CLKOUT0; // @[Buf.scala 34:26]
  assign apb0Pclk_pad_1_I = apb0Pclk_pad_O; // @[HBMDriver.scala 63:63]
  assign apb0Pclk_pad_2_I = apb0Pclk_pad_1_O; // @[HBMDriver.scala 63:71]
  assign axiAclkIn0_pad_I = mmcmGlbl_io_CLKOUT1; // @[Buf.scala 34:26]
  assign hbmRefClk0_pad_I = mmcmGlbl_io_CLKOUT2; // @[Buf.scala 34:26]
  assign apb1Pclk_pad_I = mmcmGlbl_io_CLKOUT3; // @[Buf.scala 34:26]
  assign apb1Pclk_pad_1_I = apb1Pclk_pad_O; // @[HBMDriver.scala 66:63]
  assign apb1Pclk_pad_2_I = apb1Pclk_pad_1_O; // @[HBMDriver.scala 66:71]
  assign axiAclkIn1_pad_I = mmcmGlbl_io_CLKOUT4; // @[Buf.scala 34:26]
  assign hbmRefClk1_pad_I = mmcmGlbl_io_CLKOUT5; // @[Buf.scala 34:26]
  assign mmcmAxi_io_CLKIN1 = axiAclkIn0_pad_O; // @[HBMDriver.scala 84:33]
  assign mmcmAxi_io_RST = ~mmcmGlbl_io_LOCKED; // @[HBMDriver.scala 85:36]
  assign axiAclk_pad_I = mmcmAxi_io_CLKOUT0; // @[Buf.scala 34:26]
  assign instHbm_HBM_REF_CLK_0 = hbmRefClk0_pad_O; // @[HBMDriver.scala 103:41]
  assign instHbm_HBM_REF_CLK_1 = hbmRefClk1_pad_O; // @[HBMDriver.scala 104:41]
  assign instHbm_AXI_00_ACLK = axiAclk_pad_O; // @[HBMDriver.scala 115:49]
  assign instHbm_AXI_00_ARESET_N = mmcmAxi_io_LOCKED; // @[HBMDriver.scala 116:49]
  assign instHbm_AXI_00_ARADDR = 33'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_00_ARBURST = 2'h1; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_00_ARID = 6'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_00_ARLEN = 4'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_00_ARSIZE = 3'h5; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_00_ARVALID = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_00_AWADDR = 33'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_00_AWBURST = 2'h1; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_00_AWID = 6'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_00_AWLEN = 4'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_00_AWSIZE = 3'h5; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_00_AWVALID = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_00_WDATA = 256'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_00_WLAST = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_00_WSTRB = 32'hffffffff; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_00_WVALID = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_00_RREADY = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_00_BREADY = 1'h1; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_00_WDATA_PARITY = 32'h0; // @[HBMDriver.scala 146:49]
  assign instHbm_AXI_01_ACLK = axiAclk_pad_O; // @[HBMDriver.scala 149:49]
  assign instHbm_AXI_01_ARESET_N = mmcmAxi_io_LOCKED; // @[HBMDriver.scala 150:49]
  assign instHbm_AXI_01_ARADDR = 33'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_01_ARBURST = 2'h1; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_01_ARID = 6'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_01_ARLEN = 4'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_01_ARSIZE = 3'h5; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_01_ARVALID = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_01_AWADDR = 33'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_01_AWBURST = 2'h1; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_01_AWID = 6'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_01_AWLEN = 4'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_01_AWSIZE = 3'h5; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_01_AWVALID = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_01_WDATA = 256'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_01_WLAST = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_01_WSTRB = 32'hffffffff; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_01_WVALID = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_01_RREADY = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_01_BREADY = 1'h1; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_01_WDATA_PARITY = 32'h0; // @[HBMDriver.scala 180:49]
  assign instHbm_AXI_02_ACLK = axiAclk_pad_O; // @[HBMDriver.scala 183:49]
  assign instHbm_AXI_02_ARESET_N = mmcmAxi_io_LOCKED; // @[HBMDriver.scala 184:49]
  assign instHbm_AXI_02_ARADDR = 33'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_02_ARBURST = 2'h1; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_02_ARID = 6'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_02_ARLEN = 4'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_02_ARSIZE = 3'h5; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_02_ARVALID = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_02_AWADDR = 33'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_02_AWBURST = 2'h1; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_02_AWID = 6'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_02_AWLEN = 4'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_02_AWSIZE = 3'h5; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_02_AWVALID = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_02_WDATA = 256'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_02_WLAST = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_02_WSTRB = 32'hffffffff; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_02_WVALID = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_02_RREADY = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_02_BREADY = 1'h1; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_02_WDATA_PARITY = 32'h0; // @[HBMDriver.scala 214:49]
  assign instHbm_AXI_03_ACLK = axiAclk_pad_O; // @[HBMDriver.scala 217:49]
  assign instHbm_AXI_03_ARESET_N = mmcmAxi_io_LOCKED; // @[HBMDriver.scala 218:49]
  assign instHbm_AXI_03_ARADDR = 33'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_03_ARBURST = 2'h1; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_03_ARID = 6'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_03_ARLEN = 4'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_03_ARSIZE = 3'h5; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_03_ARVALID = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_03_AWADDR = 33'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_03_AWBURST = 2'h1; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_03_AWID = 6'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_03_AWLEN = 4'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_03_AWSIZE = 3'h5; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_03_AWVALID = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_03_WDATA = 256'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_03_WLAST = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_03_WSTRB = 32'hffffffff; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_03_WVALID = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_03_RREADY = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_03_BREADY = 1'h1; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_03_WDATA_PARITY = 32'h0; // @[HBMDriver.scala 248:49]
  assign instHbm_AXI_04_ACLK = axiAclk_pad_O; // @[HBMDriver.scala 251:49]
  assign instHbm_AXI_04_ARESET_N = mmcmAxi_io_LOCKED; // @[HBMDriver.scala 252:49]
  assign instHbm_AXI_04_ARADDR = 33'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_04_ARBURST = 2'h1; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_04_ARID = 6'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_04_ARLEN = 4'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_04_ARSIZE = 3'h5; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_04_ARVALID = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_04_AWADDR = 33'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_04_AWBURST = 2'h1; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_04_AWID = 6'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_04_AWLEN = 4'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_04_AWSIZE = 3'h5; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_04_AWVALID = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_04_WDATA = 256'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_04_WLAST = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_04_WSTRB = 32'hffffffff; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_04_WVALID = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_04_RREADY = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_04_BREADY = 1'h1; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_04_WDATA_PARITY = 32'h0; // @[HBMDriver.scala 282:49]
  assign instHbm_AXI_05_ACLK = axiAclk_pad_O; // @[HBMDriver.scala 285:49]
  assign instHbm_AXI_05_ARESET_N = mmcmAxi_io_LOCKED; // @[HBMDriver.scala 286:49]
  assign instHbm_AXI_05_ARADDR = 33'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_05_ARBURST = 2'h1; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_05_ARID = 6'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_05_ARLEN = 4'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_05_ARSIZE = 3'h5; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_05_ARVALID = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_05_AWADDR = 33'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_05_AWBURST = 2'h1; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_05_AWID = 6'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_05_AWLEN = 4'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_05_AWSIZE = 3'h5; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_05_AWVALID = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_05_WDATA = 256'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_05_WLAST = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_05_WSTRB = 32'hffffffff; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_05_WVALID = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_05_RREADY = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_05_BREADY = 1'h1; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_05_WDATA_PARITY = 32'h0; // @[HBMDriver.scala 316:49]
  assign instHbm_AXI_06_ACLK = axiAclk_pad_O; // @[HBMDriver.scala 319:49]
  assign instHbm_AXI_06_ARESET_N = mmcmAxi_io_LOCKED; // @[HBMDriver.scala 320:49]
  assign instHbm_AXI_06_ARADDR = 33'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_06_ARBURST = 2'h1; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_06_ARID = 6'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_06_ARLEN = 4'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_06_ARSIZE = 3'h5; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_06_ARVALID = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_06_AWADDR = 33'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_06_AWBURST = 2'h1; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_06_AWID = 6'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_06_AWLEN = 4'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_06_AWSIZE = 3'h5; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_06_AWVALID = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_06_WDATA = 256'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_06_WLAST = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_06_WSTRB = 32'hffffffff; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_06_WVALID = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_06_RREADY = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_06_BREADY = 1'h1; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_06_WDATA_PARITY = 32'h0; // @[HBMDriver.scala 350:49]
  assign instHbm_AXI_07_ACLK = axiAclk_pad_O; // @[HBMDriver.scala 353:49]
  assign instHbm_AXI_07_ARESET_N = mmcmAxi_io_LOCKED; // @[HBMDriver.scala 354:49]
  assign instHbm_AXI_07_ARADDR = 33'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_07_ARBURST = 2'h1; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_07_ARID = 6'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_07_ARLEN = 4'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_07_ARSIZE = 3'h5; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_07_ARVALID = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_07_AWADDR = 33'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_07_AWBURST = 2'h1; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_07_AWID = 6'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_07_AWLEN = 4'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_07_AWSIZE = 3'h5; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_07_AWVALID = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_07_WDATA = 256'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_07_WLAST = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_07_WSTRB = 32'hffffffff; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_07_WVALID = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_07_RREADY = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_07_BREADY = 1'h1; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_07_WDATA_PARITY = 32'h0; // @[HBMDriver.scala 384:49]
  assign instHbm_AXI_08_ACLK = axiAclk_pad_O; // @[HBMDriver.scala 387:49]
  assign instHbm_AXI_08_ARESET_N = mmcmAxi_io_LOCKED; // @[HBMDriver.scala 388:49]
  assign instHbm_AXI_08_ARADDR = 33'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_08_ARBURST = 2'h1; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_08_ARID = 6'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_08_ARLEN = 4'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_08_ARSIZE = 3'h5; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_08_ARVALID = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_08_AWADDR = 33'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_08_AWBURST = 2'h1; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_08_AWID = 6'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_08_AWLEN = 4'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_08_AWSIZE = 3'h5; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_08_AWVALID = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_08_WDATA = 256'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_08_WLAST = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_08_WSTRB = 32'hffffffff; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_08_WVALID = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_08_RREADY = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_08_BREADY = 1'h1; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_08_WDATA_PARITY = 32'h0; // @[HBMDriver.scala 418:49]
  assign instHbm_AXI_09_ACLK = axiAclk_pad_O; // @[HBMDriver.scala 421:49]
  assign instHbm_AXI_09_ARESET_N = mmcmAxi_io_LOCKED; // @[HBMDriver.scala 422:49]
  assign instHbm_AXI_09_ARADDR = 33'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_09_ARBURST = 2'h1; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_09_ARID = 6'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_09_ARLEN = 4'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_09_ARSIZE = 3'h5; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_09_ARVALID = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_09_AWADDR = 33'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_09_AWBURST = 2'h1; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_09_AWID = 6'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_09_AWLEN = 4'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_09_AWSIZE = 3'h5; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_09_AWVALID = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_09_WDATA = 256'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_09_WLAST = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_09_WSTRB = 32'hffffffff; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_09_WVALID = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_09_RREADY = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_09_BREADY = 1'h1; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_09_WDATA_PARITY = 32'h0; // @[HBMDriver.scala 452:49]
  assign instHbm_AXI_10_ACLK = axiAclk_pad_O; // @[HBMDriver.scala 455:49]
  assign instHbm_AXI_10_ARESET_N = mmcmAxi_io_LOCKED; // @[HBMDriver.scala 456:49]
  assign instHbm_AXI_10_ARADDR = 33'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_10_ARBURST = 2'h1; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_10_ARID = 6'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_10_ARLEN = 4'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_10_ARSIZE = 3'h5; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_10_ARVALID = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_10_AWADDR = 33'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_10_AWBURST = 2'h1; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_10_AWID = 6'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_10_AWLEN = 4'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_10_AWSIZE = 3'h5; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_10_AWVALID = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_10_WDATA = 256'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_10_WLAST = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_10_WSTRB = 32'hffffffff; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_10_WVALID = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_10_RREADY = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_10_BREADY = 1'h1; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_10_WDATA_PARITY = 32'h0; // @[HBMDriver.scala 486:49]
  assign instHbm_AXI_11_ACLK = axiAclk_pad_O; // @[HBMDriver.scala 489:49]
  assign instHbm_AXI_11_ARESET_N = mmcmAxi_io_LOCKED; // @[HBMDriver.scala 490:49]
  assign instHbm_AXI_11_ARADDR = 33'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_11_ARBURST = 2'h1; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_11_ARID = 6'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_11_ARLEN = 4'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_11_ARSIZE = 3'h5; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_11_ARVALID = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_11_AWADDR = 33'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_11_AWBURST = 2'h1; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_11_AWID = 6'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_11_AWLEN = 4'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_11_AWSIZE = 3'h5; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_11_AWVALID = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_11_WDATA = 256'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_11_WLAST = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_11_WSTRB = 32'hffffffff; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_11_WVALID = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_11_RREADY = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_11_BREADY = 1'h1; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_11_WDATA_PARITY = 32'h0; // @[HBMDriver.scala 520:49]
  assign instHbm_AXI_12_ACLK = axiAclk_pad_O; // @[HBMDriver.scala 523:49]
  assign instHbm_AXI_12_ARESET_N = mmcmAxi_io_LOCKED; // @[HBMDriver.scala 524:49]
  assign instHbm_AXI_12_ARADDR = 33'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_12_ARBURST = 2'h1; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_12_ARID = 6'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_12_ARLEN = 4'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_12_ARSIZE = 3'h5; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_12_ARVALID = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_12_AWADDR = 33'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_12_AWBURST = 2'h1; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_12_AWID = 6'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_12_AWLEN = 4'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_12_AWSIZE = 3'h5; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_12_AWVALID = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_12_WDATA = 256'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_12_WLAST = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_12_WSTRB = 32'hffffffff; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_12_WVALID = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_12_RREADY = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_12_BREADY = 1'h1; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_12_WDATA_PARITY = 32'h0; // @[HBMDriver.scala 554:49]
  assign instHbm_AXI_13_ACLK = axiAclk_pad_O; // @[HBMDriver.scala 557:49]
  assign instHbm_AXI_13_ARESET_N = mmcmAxi_io_LOCKED; // @[HBMDriver.scala 558:49]
  assign instHbm_AXI_13_ARADDR = 33'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_13_ARBURST = 2'h1; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_13_ARID = 6'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_13_ARLEN = 4'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_13_ARSIZE = 3'h5; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_13_ARVALID = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_13_AWADDR = 33'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_13_AWBURST = 2'h1; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_13_AWID = 6'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_13_AWLEN = 4'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_13_AWSIZE = 3'h5; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_13_AWVALID = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_13_WDATA = 256'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_13_WLAST = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_13_WSTRB = 32'hffffffff; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_13_WVALID = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_13_RREADY = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_13_BREADY = 1'h1; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_13_WDATA_PARITY = 32'h0; // @[HBMDriver.scala 588:49]
  assign instHbm_AXI_14_ACLK = axiAclk_pad_O; // @[HBMDriver.scala 591:49]
  assign instHbm_AXI_14_ARESET_N = mmcmAxi_io_LOCKED; // @[HBMDriver.scala 592:49]
  assign instHbm_AXI_14_ARADDR = 33'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_14_ARBURST = 2'h1; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_14_ARID = 6'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_14_ARLEN = 4'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_14_ARSIZE = 3'h5; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_14_ARVALID = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_14_AWADDR = 33'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_14_AWBURST = 2'h1; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_14_AWID = 6'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_14_AWLEN = 4'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_14_AWSIZE = 3'h5; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_14_AWVALID = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_14_WDATA = 256'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_14_WLAST = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_14_WSTRB = 32'hffffffff; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_14_WVALID = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_14_RREADY = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_14_BREADY = 1'h1; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_14_WDATA_PARITY = 32'h0; // @[HBMDriver.scala 622:49]
  assign instHbm_AXI_15_ACLK = axiAclk_pad_O; // @[HBMDriver.scala 625:49]
  assign instHbm_AXI_15_ARESET_N = mmcmAxi_io_LOCKED; // @[HBMDriver.scala 626:49]
  assign instHbm_AXI_15_ARADDR = 33'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_15_ARBURST = 2'h1; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_15_ARID = 6'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_15_ARLEN = 4'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_15_ARSIZE = 3'h5; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_15_ARVALID = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_15_AWADDR = 33'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_15_AWBURST = 2'h1; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_15_AWID = 6'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_15_AWLEN = 4'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_15_AWSIZE = 3'h5; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_15_AWVALID = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_15_WDATA = 256'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_15_WLAST = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_15_WSTRB = 32'hffffffff; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_15_WVALID = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_15_RREADY = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_15_BREADY = 1'h1; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_15_WDATA_PARITY = 32'h0; // @[HBMDriver.scala 656:49]
  assign instHbm_AXI_16_ACLK = axiAclk_pad_O; // @[HBMDriver.scala 667:49]
  assign instHbm_AXI_16_ARESET_N = mmcmAxi_io_LOCKED; // @[HBMDriver.scala 668:49]
  assign instHbm_AXI_16_ARADDR = 33'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_16_ARBURST = 2'h1; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_16_ARID = 6'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_16_ARLEN = 4'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_16_ARSIZE = 3'h5; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_16_ARVALID = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_16_AWADDR = 33'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_16_AWBURST = 2'h1; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_16_AWID = 6'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_16_AWLEN = 4'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_16_AWSIZE = 3'h5; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_16_AWVALID = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_16_WDATA = 256'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_16_WLAST = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_16_WSTRB = 32'hffffffff; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_16_WVALID = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_16_RREADY = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_16_BREADY = 1'h1; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_16_WDATA_PARITY = 32'h0; // @[HBMDriver.scala 698:49]
  assign instHbm_AXI_17_ACLK = axiAclk_pad_O; // @[HBMDriver.scala 701:49]
  assign instHbm_AXI_17_ARESET_N = mmcmAxi_io_LOCKED; // @[HBMDriver.scala 702:49]
  assign instHbm_AXI_17_ARADDR = 33'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_17_ARBURST = 2'h1; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_17_ARID = 6'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_17_ARLEN = 4'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_17_ARSIZE = 3'h5; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_17_ARVALID = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_17_AWADDR = 33'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_17_AWBURST = 2'h1; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_17_AWID = 6'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_17_AWLEN = 4'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_17_AWSIZE = 3'h5; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_17_AWVALID = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_17_WDATA = 256'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_17_WLAST = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_17_WSTRB = 32'hffffffff; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_17_WVALID = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_17_RREADY = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_17_BREADY = 1'h1; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_17_WDATA_PARITY = 32'h0; // @[HBMDriver.scala 732:49]
  assign instHbm_AXI_18_ACLK = axiAclk_pad_O; // @[HBMDriver.scala 735:49]
  assign instHbm_AXI_18_ARESET_N = mmcmAxi_io_LOCKED; // @[HBMDriver.scala 736:49]
  assign instHbm_AXI_18_ARADDR = 33'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_18_ARBURST = 2'h1; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_18_ARID = 6'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_18_ARLEN = 4'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_18_ARSIZE = 3'h5; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_18_ARVALID = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_18_AWADDR = 33'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_18_AWBURST = 2'h1; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_18_AWID = 6'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_18_AWLEN = 4'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_18_AWSIZE = 3'h5; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_18_AWVALID = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_18_WDATA = 256'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_18_WLAST = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_18_WSTRB = 32'hffffffff; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_18_WVALID = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_18_RREADY = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_18_BREADY = 1'h1; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_18_WDATA_PARITY = 32'h0; // @[HBMDriver.scala 766:49]
  assign instHbm_AXI_19_ACLK = axiAclk_pad_O; // @[HBMDriver.scala 769:49]
  assign instHbm_AXI_19_ARESET_N = mmcmAxi_io_LOCKED; // @[HBMDriver.scala 770:49]
  assign instHbm_AXI_19_ARADDR = 33'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_19_ARBURST = 2'h1; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_19_ARID = 6'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_19_ARLEN = 4'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_19_ARSIZE = 3'h5; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_19_ARVALID = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_19_AWADDR = 33'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_19_AWBURST = 2'h1; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_19_AWID = 6'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_19_AWLEN = 4'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_19_AWSIZE = 3'h5; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_19_AWVALID = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_19_WDATA = 256'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_19_WLAST = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_19_WSTRB = 32'hffffffff; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_19_WVALID = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_19_RREADY = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_19_BREADY = 1'h1; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_19_WDATA_PARITY = 32'h0; // @[HBMDriver.scala 800:49]
  assign instHbm_AXI_20_ACLK = axiAclk_pad_O; // @[HBMDriver.scala 803:49]
  assign instHbm_AXI_20_ARESET_N = mmcmAxi_io_LOCKED; // @[HBMDriver.scala 804:49]
  assign instHbm_AXI_20_ARADDR = 33'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_20_ARBURST = 2'h1; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_20_ARID = 6'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_20_ARLEN = 4'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_20_ARSIZE = 3'h5; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_20_ARVALID = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_20_AWADDR = 33'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_20_AWBURST = 2'h1; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_20_AWID = 6'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_20_AWLEN = 4'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_20_AWSIZE = 3'h5; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_20_AWVALID = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_20_WDATA = 256'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_20_WLAST = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_20_WSTRB = 32'hffffffff; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_20_WVALID = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_20_RREADY = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_20_BREADY = 1'h1; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_20_WDATA_PARITY = 32'h0; // @[HBMDriver.scala 834:49]
  assign instHbm_AXI_21_ACLK = axiAclk_pad_O; // @[HBMDriver.scala 837:49]
  assign instHbm_AXI_21_ARESET_N = mmcmAxi_io_LOCKED; // @[HBMDriver.scala 838:49]
  assign instHbm_AXI_21_ARADDR = 33'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_21_ARBURST = 2'h1; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_21_ARID = 6'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_21_ARLEN = 4'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_21_ARSIZE = 3'h5; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_21_ARVALID = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_21_AWADDR = 33'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_21_AWBURST = 2'h1; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_21_AWID = 6'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_21_AWLEN = 4'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_21_AWSIZE = 3'h5; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_21_AWVALID = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_21_WDATA = 256'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_21_WLAST = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_21_WSTRB = 32'hffffffff; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_21_WVALID = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_21_RREADY = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_21_BREADY = 1'h1; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_21_WDATA_PARITY = 32'h0; // @[HBMDriver.scala 868:49]
  assign instHbm_AXI_22_ACLK = axiAclk_pad_O; // @[HBMDriver.scala 871:49]
  assign instHbm_AXI_22_ARESET_N = mmcmAxi_io_LOCKED; // @[HBMDriver.scala 872:49]
  assign instHbm_AXI_22_ARADDR = 33'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_22_ARBURST = 2'h1; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_22_ARID = 6'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_22_ARLEN = 4'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_22_ARSIZE = 3'h5; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_22_ARVALID = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_22_AWADDR = 33'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_22_AWBURST = 2'h1; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_22_AWID = 6'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_22_AWLEN = 4'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_22_AWSIZE = 3'h5; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_22_AWVALID = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_22_WDATA = 256'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_22_WLAST = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_22_WSTRB = 32'hffffffff; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_22_WVALID = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_22_RREADY = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_22_BREADY = 1'h1; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_22_WDATA_PARITY = 32'h0; // @[HBMDriver.scala 902:49]
  assign instHbm_AXI_23_ACLK = axiAclk_pad_O; // @[HBMDriver.scala 905:49]
  assign instHbm_AXI_23_ARESET_N = mmcmAxi_io_LOCKED; // @[HBMDriver.scala 906:49]
  assign instHbm_AXI_23_ARADDR = 33'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_23_ARBURST = 2'h1; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_23_ARID = 6'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_23_ARLEN = 4'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_23_ARSIZE = 3'h5; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_23_ARVALID = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_23_AWADDR = 33'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_23_AWBURST = 2'h1; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_23_AWID = 6'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_23_AWLEN = 4'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_23_AWSIZE = 3'h5; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_23_AWVALID = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_23_WDATA = 256'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_23_WLAST = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_23_WSTRB = 32'hffffffff; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_23_WVALID = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_23_RREADY = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_23_BREADY = 1'h1; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_23_WDATA_PARITY = 32'h0; // @[HBMDriver.scala 936:49]
  assign instHbm_AXI_24_ACLK = axiAclk_pad_O; // @[HBMDriver.scala 939:49]
  assign instHbm_AXI_24_ARESET_N = mmcmAxi_io_LOCKED; // @[HBMDriver.scala 940:49]
  assign instHbm_AXI_24_ARADDR = 33'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_24_ARBURST = 2'h1; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_24_ARID = 6'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_24_ARLEN = 4'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_24_ARSIZE = 3'h5; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_24_ARVALID = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_24_AWADDR = 33'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_24_AWBURST = 2'h1; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_24_AWID = 6'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_24_AWLEN = 4'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_24_AWSIZE = 3'h5; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_24_AWVALID = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_24_WDATA = 256'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_24_WLAST = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_24_WSTRB = 32'hffffffff; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_24_WVALID = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_24_RREADY = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_24_BREADY = 1'h1; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_24_WDATA_PARITY = 32'h0; // @[HBMDriver.scala 970:49]
  assign instHbm_AXI_25_ACLK = axiAclk_pad_O; // @[HBMDriver.scala 973:49]
  assign instHbm_AXI_25_ARESET_N = mmcmAxi_io_LOCKED; // @[HBMDriver.scala 974:49]
  assign instHbm_AXI_25_ARADDR = 33'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_25_ARBURST = 2'h1; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_25_ARID = 6'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_25_ARLEN = 4'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_25_ARSIZE = 3'h5; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_25_ARVALID = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_25_AWADDR = 33'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_25_AWBURST = 2'h1; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_25_AWID = 6'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_25_AWLEN = 4'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_25_AWSIZE = 3'h5; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_25_AWVALID = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_25_WDATA = 256'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_25_WLAST = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_25_WSTRB = 32'hffffffff; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_25_WVALID = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_25_RREADY = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_25_BREADY = 1'h1; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_25_WDATA_PARITY = 32'h0; // @[HBMDriver.scala 1004:49]
  assign instHbm_AXI_26_ACLK = axiAclk_pad_O; // @[HBMDriver.scala 1007:49]
  assign instHbm_AXI_26_ARESET_N = mmcmAxi_io_LOCKED; // @[HBMDriver.scala 1008:49]
  assign instHbm_AXI_26_ARADDR = 33'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_26_ARBURST = 2'h1; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_26_ARID = 6'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_26_ARLEN = 4'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_26_ARSIZE = 3'h5; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_26_ARVALID = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_26_AWADDR = 33'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_26_AWBURST = 2'h1; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_26_AWID = 6'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_26_AWLEN = 4'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_26_AWSIZE = 3'h5; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_26_AWVALID = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_26_WDATA = 256'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_26_WLAST = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_26_WSTRB = 32'hffffffff; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_26_WVALID = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_26_RREADY = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_26_BREADY = 1'h1; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_26_WDATA_PARITY = 32'h0; // @[HBMDriver.scala 1038:49]
  assign instHbm_AXI_27_ACLK = axiAclk_pad_O; // @[HBMDriver.scala 1041:49]
  assign instHbm_AXI_27_ARESET_N = mmcmAxi_io_LOCKED; // @[HBMDriver.scala 1042:49]
  assign instHbm_AXI_27_ARADDR = 33'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_27_ARBURST = 2'h1; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_27_ARID = 6'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_27_ARLEN = 4'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_27_ARSIZE = 3'h5; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_27_ARVALID = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_27_AWADDR = 33'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_27_AWBURST = 2'h1; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_27_AWID = 6'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_27_AWLEN = 4'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_27_AWSIZE = 3'h5; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_27_AWVALID = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_27_WDATA = 256'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_27_WLAST = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_27_WSTRB = 32'hffffffff; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_27_WVALID = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_27_RREADY = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_27_BREADY = 1'h1; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_27_WDATA_PARITY = 32'h0; // @[HBMDriver.scala 1072:49]
  assign instHbm_AXI_28_ACLK = axiAclk_pad_O; // @[HBMDriver.scala 1075:49]
  assign instHbm_AXI_28_ARESET_N = mmcmAxi_io_LOCKED; // @[HBMDriver.scala 1076:49]
  assign instHbm_AXI_28_ARADDR = 33'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_28_ARBURST = 2'h1; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_28_ARID = 6'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_28_ARLEN = 4'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_28_ARSIZE = 3'h5; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_28_ARVALID = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_28_AWADDR = 33'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_28_AWBURST = 2'h1; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_28_AWID = 6'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_28_AWLEN = 4'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_28_AWSIZE = 3'h5; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_28_AWVALID = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_28_WDATA = 256'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_28_WLAST = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_28_WSTRB = 32'hffffffff; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_28_WVALID = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_28_RREADY = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_28_BREADY = 1'h1; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_28_WDATA_PARITY = 32'h0; // @[HBMDriver.scala 1106:49]
  assign instHbm_AXI_29_ACLK = axiAclk_pad_O; // @[HBMDriver.scala 1109:49]
  assign instHbm_AXI_29_ARESET_N = mmcmAxi_io_LOCKED; // @[HBMDriver.scala 1110:49]
  assign instHbm_AXI_29_ARADDR = 33'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_29_ARBURST = 2'h1; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_29_ARID = 6'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_29_ARLEN = 4'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_29_ARSIZE = 3'h5; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_29_ARVALID = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_29_AWADDR = 33'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_29_AWBURST = 2'h1; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_29_AWID = 6'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_29_AWLEN = 4'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_29_AWSIZE = 3'h5; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_29_AWVALID = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_29_WDATA = 256'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_29_WLAST = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_29_WSTRB = 32'hffffffff; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_29_WVALID = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_29_RREADY = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_29_BREADY = 1'h1; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_29_WDATA_PARITY = 32'h0; // @[HBMDriver.scala 1140:49]
  assign instHbm_AXI_30_ACLK = axiAclk_pad_O; // @[HBMDriver.scala 1143:49]
  assign instHbm_AXI_30_ARESET_N = mmcmAxi_io_LOCKED; // @[HBMDriver.scala 1144:49]
  assign instHbm_AXI_30_ARADDR = 33'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_30_ARBURST = 2'h1; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_30_ARID = 6'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_30_ARLEN = 4'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_30_ARSIZE = 3'h5; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_30_ARVALID = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_30_AWADDR = 33'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_30_AWBURST = 2'h1; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_30_AWID = 6'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_30_AWLEN = 4'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_30_AWSIZE = 3'h5; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_30_AWVALID = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_30_WDATA = 256'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_30_WLAST = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_30_WSTRB = 32'hffffffff; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_30_WVALID = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_30_RREADY = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_30_BREADY = 1'h1; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_30_WDATA_PARITY = 32'h0; // @[HBMDriver.scala 1174:49]
  assign instHbm_AXI_31_ACLK = axiAclk_pad_O; // @[HBMDriver.scala 1177:49]
  assign instHbm_AXI_31_ARESET_N = mmcmAxi_io_LOCKED; // @[HBMDriver.scala 1178:49]
  assign instHbm_AXI_31_ARADDR = 33'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_31_ARBURST = 2'h1; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_31_ARID = 6'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_31_ARLEN = 4'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_31_ARSIZE = 3'h5; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_31_ARVALID = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_31_AWADDR = 33'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_31_AWBURST = 2'h1; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_31_AWID = 6'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_31_AWLEN = 4'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_31_AWSIZE = 3'h5; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_31_AWVALID = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_31_WDATA = 256'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_31_WLAST = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_31_WSTRB = 32'hffffffff; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_31_WVALID = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_31_RREADY = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_31_BREADY = 1'h1; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_31_WDATA_PARITY = 32'h0; // @[HBMDriver.scala 1208:49]
  assign instHbm_APB_0_PWDATA = 32'h0; // @[HBMDriver.scala 1214:36]
  assign instHbm_APB_0_PADDR = 22'h0; // @[HBMDriver.scala 1215:36]
  assign instHbm_APB_0_PCLK = apb0Pclk_pad_2_O; // @[HBMDriver.scala 1216:36]
  assign instHbm_APB_0_PENABLE = 1'h0; // @[HBMDriver.scala 1217:36]
  assign instHbm_APB_0_PRESET_N = mmcmGlbl_io_LOCKED; // @[HBMDriver.scala 1218:36]
  assign instHbm_APB_0_PSEL = 1'h0; // @[HBMDriver.scala 1219:36]
  assign instHbm_APB_0_PWRITE = 1'h0; // @[HBMDriver.scala 1220:36]
  assign instHbm_APB_1_PWDATA = 32'h0; // @[HBMDriver.scala 1225:36]
  assign instHbm_APB_1_PADDR = 22'h0; // @[HBMDriver.scala 1226:36]
  assign instHbm_APB_1_PCLK = apb1Pclk_pad_2_O; // @[HBMDriver.scala 1227:36]
  assign instHbm_APB_1_PENABLE = 1'h0; // @[HBMDriver.scala 1228:36]
  assign instHbm_APB_1_PRESET_N = mmcmGlbl_io_LOCKED; // @[HBMDriver.scala 1229:36]
  assign instHbm_APB_1_PSEL = 1'h0; // @[HBMDriver.scala 1230:36]
  assign instHbm_APB_1_PWRITE = 1'h0; // @[HBMDriver.scala 1231:36]
  always @(posedge apb0Pclk_pad_2_O) begin
    apb_complete_0_r <= instHbm_apb_complete_0; // @[Reg.scala 16:19 Reg.scala 16:23 Reg.scala 15:16]
    apb_complete_0 <= apb_complete_0_r; // @[Reg.scala 16:19 Reg.scala 16:23 Reg.scala 15:16]
  end
  always @(posedge apb1Pclk_pad_2_O) begin
    apb_complete_1_r <= instHbm_apb_complete_1; // @[Reg.scala 16:19 Reg.scala 16:23 Reg.scala 15:16]
    apb_complete_1 <= apb_complete_1_r; // @[Reg.scala 16:19 Reg.scala 16:23 Reg.scala 15:16]
  end
  always @(posedge axiAclk_pad_O) begin
    io_hbm_rstn_REG <= mmcmAxi_io_LOCKED; // @[HBMDriver.scala 97:63]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  apb_complete_0_r = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  apb_complete_0 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  apb_complete_1_r = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  apb_complete_1 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  io_hbm_rstn_REG = _RAND_4[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module SV_STREAM_FIFO(
  input          io_m_clk,
  input          io_s_clk,
  input          io_reset_n,
  input  [599:0] io_in_data,
  input          io_in_valid,
  output         io_in_ready,
  output         io_out_valid
);
  wire [599:0] meta_m_axis_tdata; // @[Meta.scala 30:26]
  wire [74:0] meta_m_axis_tkeep; // @[Meta.scala 30:26]
  wire  meta_m_axis_tlast; // @[Meta.scala 30:26]
  wire  meta_m_axis_tvalid; // @[Meta.scala 30:26]
  wire [4:0] meta_rd_data_count_axis; // @[Meta.scala 30:26]
  wire  meta_s_axis_tready; // @[Meta.scala 30:26]
  wire [4:0] meta_wr_data_count_axis; // @[Meta.scala 30:26]
  wire  meta_m_aclk; // @[Meta.scala 30:26]
  wire  meta_m_axis_tready; // @[Meta.scala 30:26]
  wire  meta_s_aclk; // @[Meta.scala 30:26]
  wire  meta_s_aresetn; // @[Meta.scala 30:26]
  wire [599:0] meta_s_axis_tdata; // @[Meta.scala 30:26]
  wire  meta_s_axis_tdest; // @[Meta.scala 30:26]
  wire  meta_s_axis_tid; // @[Meta.scala 30:26]
  wire [74:0] meta_s_axis_tkeep; // @[Meta.scala 30:26]
  wire  meta_s_axis_tlast; // @[Meta.scala 30:26]
  wire [74:0] meta_s_axis_tstrb; // @[Meta.scala 30:26]
  wire  meta_s_axis_tuser; // @[Meta.scala 30:26]
  wire  meta_s_axis_tvalid; // @[Meta.scala 30:26]
  xpm_fifo_axis
    #(.RD_DATA_COUNT_WIDTH(5), .CLOCKING_MODE("independent_clock"), .PACKET_FIFO("false"), .USE_ADV_FEATURES("0404"), .TID_WIDTH(1), .TDEST_WIDTH(1), .PROG_EMPTY_THRESH(10), .TUSER_WIDTH(1), .FIFO_DEPTH(16), .SIM_ASSERT_CHK(0), .WR_DATA_COUNT_WIDTH(5), .ECC_MODE("no_ecc"), .FIFO_MEMORY_TYPE("auto"), .PROG_FULL_THRESH(10), .TDATA_WIDTH(600), .RELATED_CLOCKS(0), .CASCADE_HEIGHT(0), .CDC_SYNC_STAGES(2))
    meta ( // @[Meta.scala 30:26]
    .m_axis_tdata(meta_m_axis_tdata),
    .m_axis_tkeep(meta_m_axis_tkeep),
    .m_axis_tlast(meta_m_axis_tlast),
    .m_axis_tvalid(meta_m_axis_tvalid),
    .rd_data_count_axis(meta_rd_data_count_axis),
    .s_axis_tready(meta_s_axis_tready),
    .wr_data_count_axis(meta_wr_data_count_axis),
    .m_aclk(meta_m_aclk),
    .m_axis_tready(meta_m_axis_tready),
    .s_aclk(meta_s_aclk),
    .s_aresetn(meta_s_aresetn),
    .s_axis_tdata(meta_s_axis_tdata),
    .s_axis_tdest(meta_s_axis_tdest),
    .s_axis_tid(meta_s_axis_tid),
    .s_axis_tkeep(meta_s_axis_tkeep),
    .s_axis_tlast(meta_s_axis_tlast),
    .s_axis_tstrb(meta_s_axis_tstrb),
    .s_axis_tuser(meta_s_axis_tuser),
    .s_axis_tvalid(meta_s_axis_tvalid)
  );
  assign io_in_ready = meta_s_axis_tready; // @[Meta.scala 34:41]
  assign io_out_valid = meta_m_axis_tvalid; // @[Meta.scala 32:41]
  assign meta_m_aclk = io_m_clk; // @[Meta.scala 37:49]
  assign meta_m_axis_tready = 1'h1; // @[Meta.scala 38:41]
  assign meta_s_aclk = io_s_clk; // @[Meta.scala 39:49]
  assign meta_s_aresetn = io_reset_n; // @[Meta.scala 40:49]
  assign meta_s_axis_tdata = io_in_data; // @[Meta.scala 41:41]
  assign meta_s_axis_tdest = 1'h0; // @[Meta.scala 42:41]
  assign meta_s_axis_tid = 1'h0; // @[Meta.scala 43:49]
  assign meta_s_axis_tkeep = 75'h7ffffffffffffffffff; // @[Bitwise.scala 72:12]
  assign meta_s_axis_tlast = 1'h1; // @[Meta.scala 45:41]
  assign meta_s_axis_tstrb = 75'h7ffffffffffffffffff; // @[Bitwise.scala 72:12]
  assign meta_s_axis_tuser = 1'h0; // @[Meta.scala 47:41]
  assign meta_s_axis_tvalid = io_in_valid; // @[Meta.scala 48:41]
endmodule
module XConverter(
  input          io__in_clk,
  input          io__out_clk,
  input          io__rstn,
  output         io__in_ready,
  input          io__in_valid,
  input  [511:0] io__in_bits_data,
  input  [31:0]  io__in_bits_tcrc,
  input  [10:0]  io__in_bits_tuser_qid,
  input  [2:0]   io__in_bits_tuser_port_id,
  input          io__in_bits_tuser_err,
  input  [31:0]  io__in_bits_tuser_mdata,
  input  [5:0]   io__in_bits_tuser_mty,
  input          io__in_bits_tuser_zero_byte,
  input          io__in_bits_last,
  output         io__out_valid,
  output         io_in_ready,
  output         io_in_valid
);
  wire  fifo_io_m_clk; // @[XConverter.scala 97:34]
  wire  fifo_io_s_clk; // @[XConverter.scala 97:34]
  wire  fifo_io_reset_n; // @[XConverter.scala 97:34]
  wire [599:0] fifo_io_in_data; // @[XConverter.scala 97:34]
  wire  fifo_io_in_valid; // @[XConverter.scala 97:34]
  wire  fifo_io_in_ready; // @[XConverter.scala 97:34]
  wire  fifo_io_out_valid; // @[XConverter.scala 97:34]
  wire [598:0] _fifo_io_in_data_T = {io__in_bits_data,io__in_bits_tcrc,io__in_bits_tuser_qid,io__in_bits_tuser_port_id,
    io__in_bits_tuser_err,io__in_bits_tuser_mdata,io__in_bits_tuser_mty,io__in_bits_tuser_zero_byte,io__in_bits_last}; // @[XConverter.scala 103:63]
  SV_STREAM_FIFO fifo ( // @[XConverter.scala 97:34]
    .io_m_clk(fifo_io_m_clk),
    .io_s_clk(fifo_io_s_clk),
    .io_reset_n(fifo_io_reset_n),
    .io_in_data(fifo_io_in_data),
    .io_in_valid(fifo_io_in_valid),
    .io_in_ready(fifo_io_in_ready),
    .io_out_valid(fifo_io_out_valid)
  );
  assign io__in_ready = fifo_io_in_ready; // @[XConverter.scala 105:41]
  assign io__out_valid = fifo_io_out_valid; // @[XConverter.scala 108:41]
  assign io_in_ready = io__in_ready;
  assign io_in_valid = io__in_valid;
  assign fifo_io_m_clk = io__out_clk; // @[XConverter.scala 100:41]
  assign fifo_io_s_clk = io__in_clk; // @[XConverter.scala 99:41]
  assign fifo_io_reset_n = io__rstn; // @[XConverter.scala 101:41]
  assign fifo_io_in_data = {{1'd0}, _fifo_io_in_data_T}; // @[XConverter.scala 103:63]
  assign fifo_io_in_valid = io__in_valid; // @[XConverter.scala 104:41]
endmodule
module RegSlice(
  input          clock,
  input          reset,
  output         io_upStream_ready,
  input          io_upStream_valid,
  input  [511:0] io_upStream_bits_data,
  input  [31:0]  io_upStream_bits_tcrc,
  input  [10:0]  io_upStream_bits_tuser_qid,
  input  [2:0]   io_upStream_bits_tuser_port_id,
  input          io_upStream_bits_tuser_err,
  input  [31:0]  io_upStream_bits_tuser_mdata,
  input  [5:0]   io_upStream_bits_tuser_mty,
  input          io_upStream_bits_tuser_zero_byte,
  input          io_upStream_bits_last,
  input          io_downStream_ready,
  output         io_downStream_valid,
  output [511:0] io_downStream_bits_data,
  output [31:0]  io_downStream_bits_tcrc,
  output [10:0]  io_downStream_bits_tuser_qid,
  output [2:0]   io_downStream_bits_tuser_port_id,
  output         io_downStream_bits_tuser_err,
  output [31:0]  io_downStream_bits_tuser_mdata,
  output [5:0]   io_downStream_bits_tuser_mty,
  output         io_downStream_bits_tuser_zero_byte,
  output         io_downStream_bits_last
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [511:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [511:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
`endif // RANDOMIZE_REG_INIT
  reg  fwd_valid; // @[RegSlices.scala 112:34]
  reg [511:0] fwd_data_data; // @[RegSlices.scala 113:30]
  reg [31:0] fwd_data_tcrc; // @[RegSlices.scala 113:30]
  reg [10:0] fwd_data_tuser_qid; // @[RegSlices.scala 113:30]
  reg [2:0] fwd_data_tuser_port_id; // @[RegSlices.scala 113:30]
  reg  fwd_data_tuser_err; // @[RegSlices.scala 113:30]
  reg [31:0] fwd_data_tuser_mdata; // @[RegSlices.scala 113:30]
  reg [5:0] fwd_data_tuser_mty; // @[RegSlices.scala 113:30]
  reg  fwd_data_tuser_zero_byte; // @[RegSlices.scala 113:30]
  reg  fwd_data_last; // @[RegSlices.scala 113:30]
  wire  fwd_ready_s = ~fwd_valid | io_downStream_ready; // @[RegSlices.scala 115:35]
  reg  bwd_ready; // @[RegSlices.scala 123:34]
  reg [511:0] bwd_data_data; // @[RegSlices.scala 124:30]
  reg [31:0] bwd_data_tcrc; // @[RegSlices.scala 124:30]
  reg [10:0] bwd_data_tuser_qid; // @[RegSlices.scala 124:30]
  reg [2:0] bwd_data_tuser_port_id; // @[RegSlices.scala 124:30]
  reg  bwd_data_tuser_err; // @[RegSlices.scala 124:30]
  reg [31:0] bwd_data_tuser_mdata; // @[RegSlices.scala 124:30]
  reg [5:0] bwd_data_tuser_mty; // @[RegSlices.scala 124:30]
  reg  bwd_data_tuser_zero_byte; // @[RegSlices.scala 124:30]
  reg  bwd_data_last; // @[RegSlices.scala 124:30]
  wire  _fwd_valid_T = io_downStream_ready ? 1'h0 : fwd_valid; // @[RegSlices.scala 121:53]
  wire  bwd_valid_s = ~bwd_ready | io_upStream_valid; // @[RegSlices.scala 126:39]
  wire  _bwd_ready_T = io_upStream_valid ? 1'h0 : bwd_ready; // @[RegSlices.scala 132:53]
  assign io_upStream_ready = bwd_ready; // @[RegSlices.scala 107:31 RegSlices.scala 128:25]
  assign io_downStream_valid = fwd_valid; // @[RegSlices.scala 109:31 RegSlices.scala 116:21]
  assign io_downStream_bits_data = fwd_data_data; // @[RegSlices.scala 108:31 RegSlices.scala 117:25]
  assign io_downStream_bits_tcrc = fwd_data_tcrc; // @[RegSlices.scala 108:31 RegSlices.scala 117:25]
  assign io_downStream_bits_tuser_qid = fwd_data_tuser_qid; // @[RegSlices.scala 108:31 RegSlices.scala 117:25]
  assign io_downStream_bits_tuser_port_id = fwd_data_tuser_port_id; // @[RegSlices.scala 108:31 RegSlices.scala 117:25]
  assign io_downStream_bits_tuser_err = fwd_data_tuser_err; // @[RegSlices.scala 108:31 RegSlices.scala 117:25]
  assign io_downStream_bits_tuser_mdata = fwd_data_tuser_mdata; // @[RegSlices.scala 108:31 RegSlices.scala 117:25]
  assign io_downStream_bits_tuser_mty = fwd_data_tuser_mty; // @[RegSlices.scala 108:31 RegSlices.scala 117:25]
  assign io_downStream_bits_tuser_zero_byte = fwd_data_tuser_zero_byte; // @[RegSlices.scala 108:31 RegSlices.scala 117:25]
  assign io_downStream_bits_last = fwd_data_last; // @[RegSlices.scala 108:31 RegSlices.scala 117:25]
  always @(posedge clock) begin
    if (reset) begin // @[RegSlices.scala 112:34]
      fwd_valid <= 1'h0; // @[RegSlices.scala 112:34]
    end else begin
      fwd_valid <= bwd_valid_s | _fwd_valid_T; // @[RegSlices.scala 121:25]
    end
    if (fwd_ready_s) begin // @[RegSlices.scala 119:31]
      if (bwd_ready) begin // @[RegSlices.scala 127:31]
        fwd_data_data <= io_upStream_bits_data;
      end else begin
        fwd_data_data <= bwd_data_data;
      end
    end
    if (fwd_ready_s) begin // @[RegSlices.scala 119:31]
      if (bwd_ready) begin // @[RegSlices.scala 127:31]
        fwd_data_tcrc <= io_upStream_bits_tcrc;
      end else begin
        fwd_data_tcrc <= bwd_data_tcrc;
      end
    end
    if (fwd_ready_s) begin // @[RegSlices.scala 119:31]
      if (bwd_ready) begin // @[RegSlices.scala 127:31]
        fwd_data_tuser_qid <= io_upStream_bits_tuser_qid;
      end else begin
        fwd_data_tuser_qid <= bwd_data_tuser_qid;
      end
    end
    if (fwd_ready_s) begin // @[RegSlices.scala 119:31]
      if (bwd_ready) begin // @[RegSlices.scala 127:31]
        fwd_data_tuser_port_id <= io_upStream_bits_tuser_port_id;
      end else begin
        fwd_data_tuser_port_id <= bwd_data_tuser_port_id;
      end
    end
    if (fwd_ready_s) begin // @[RegSlices.scala 119:31]
      if (bwd_ready) begin // @[RegSlices.scala 127:31]
        fwd_data_tuser_err <= io_upStream_bits_tuser_err;
      end else begin
        fwd_data_tuser_err <= bwd_data_tuser_err;
      end
    end
    if (fwd_ready_s) begin // @[RegSlices.scala 119:31]
      if (bwd_ready) begin // @[RegSlices.scala 127:31]
        fwd_data_tuser_mdata <= io_upStream_bits_tuser_mdata;
      end else begin
        fwd_data_tuser_mdata <= bwd_data_tuser_mdata;
      end
    end
    if (fwd_ready_s) begin // @[RegSlices.scala 119:31]
      if (bwd_ready) begin // @[RegSlices.scala 127:31]
        fwd_data_tuser_mty <= io_upStream_bits_tuser_mty;
      end else begin
        fwd_data_tuser_mty <= bwd_data_tuser_mty;
      end
    end
    if (fwd_ready_s) begin // @[RegSlices.scala 119:31]
      if (bwd_ready) begin // @[RegSlices.scala 127:31]
        fwd_data_tuser_zero_byte <= io_upStream_bits_tuser_zero_byte;
      end else begin
        fwd_data_tuser_zero_byte <= bwd_data_tuser_zero_byte;
      end
    end
    if (fwd_ready_s) begin // @[RegSlices.scala 119:31]
      if (bwd_ready) begin // @[RegSlices.scala 127:31]
        fwd_data_last <= io_upStream_bits_last;
      end else begin
        fwd_data_last <= bwd_data_last;
      end
    end
    bwd_ready <= reset | (fwd_ready_s | _bwd_ready_T); // @[RegSlices.scala 123:34 RegSlices.scala 123:34 RegSlices.scala 132:25]
    if (bwd_ready) begin // @[RegSlices.scala 130:31]
      bwd_data_data <= io_upStream_bits_data;
    end
    if (bwd_ready) begin // @[RegSlices.scala 130:31]
      bwd_data_tcrc <= io_upStream_bits_tcrc;
    end
    if (bwd_ready) begin // @[RegSlices.scala 130:31]
      bwd_data_tuser_qid <= io_upStream_bits_tuser_qid;
    end
    if (bwd_ready) begin // @[RegSlices.scala 130:31]
      bwd_data_tuser_port_id <= io_upStream_bits_tuser_port_id;
    end
    if (bwd_ready) begin // @[RegSlices.scala 130:31]
      bwd_data_tuser_err <= io_upStream_bits_tuser_err;
    end
    if (bwd_ready) begin // @[RegSlices.scala 130:31]
      bwd_data_tuser_mdata <= io_upStream_bits_tuser_mdata;
    end
    if (bwd_ready) begin // @[RegSlices.scala 130:31]
      bwd_data_tuser_mty <= io_upStream_bits_tuser_mty;
    end
    if (bwd_ready) begin // @[RegSlices.scala 130:31]
      bwd_data_tuser_zero_byte <= io_upStream_bits_tuser_zero_byte;
    end
    if (bwd_ready) begin // @[RegSlices.scala 130:31]
      bwd_data_last <= io_upStream_bits_last;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  fwd_valid = _RAND_0[0:0];
  _RAND_1 = {16{`RANDOM}};
  fwd_data_data = _RAND_1[511:0];
  _RAND_2 = {1{`RANDOM}};
  fwd_data_tcrc = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  fwd_data_tuser_qid = _RAND_3[10:0];
  _RAND_4 = {1{`RANDOM}};
  fwd_data_tuser_port_id = _RAND_4[2:0];
  _RAND_5 = {1{`RANDOM}};
  fwd_data_tuser_err = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  fwd_data_tuser_mdata = _RAND_6[31:0];
  _RAND_7 = {1{`RANDOM}};
  fwd_data_tuser_mty = _RAND_7[5:0];
  _RAND_8 = {1{`RANDOM}};
  fwd_data_tuser_zero_byte = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  fwd_data_last = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  bwd_ready = _RAND_10[0:0];
  _RAND_11 = {16{`RANDOM}};
  bwd_data_data = _RAND_11[511:0];
  _RAND_12 = {1{`RANDOM}};
  bwd_data_tcrc = _RAND_12[31:0];
  _RAND_13 = {1{`RANDOM}};
  bwd_data_tuser_qid = _RAND_13[10:0];
  _RAND_14 = {1{`RANDOM}};
  bwd_data_tuser_port_id = _RAND_14[2:0];
  _RAND_15 = {1{`RANDOM}};
  bwd_data_tuser_err = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  bwd_data_tuser_mdata = _RAND_16[31:0];
  _RAND_17 = {1{`RANDOM}};
  bwd_data_tuser_mty = _RAND_17[5:0];
  _RAND_18 = {1{`RANDOM}};
  bwd_data_tuser_zero_byte = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  bwd_data_last = _RAND_19[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module SV_STREAM_FIFO_1(
  input          io_m_clk,
  input          io_s_clk,
  input          io_reset_n,
  input  [607:0] io_in_data,
  input          io_in_valid,
  output         io_in_ready,
  output [607:0] io_out_data,
  output         io_out_valid,
  input          io_out_ready
);
  wire [607:0] meta_m_axis_tdata; // @[Meta.scala 30:26]
  wire [75:0] meta_m_axis_tkeep; // @[Meta.scala 30:26]
  wire  meta_m_axis_tlast; // @[Meta.scala 30:26]
  wire  meta_m_axis_tvalid; // @[Meta.scala 30:26]
  wire [4:0] meta_rd_data_count_axis; // @[Meta.scala 30:26]
  wire  meta_s_axis_tready; // @[Meta.scala 30:26]
  wire [4:0] meta_wr_data_count_axis; // @[Meta.scala 30:26]
  wire  meta_m_aclk; // @[Meta.scala 30:26]
  wire  meta_m_axis_tready; // @[Meta.scala 30:26]
  wire  meta_s_aclk; // @[Meta.scala 30:26]
  wire  meta_s_aresetn; // @[Meta.scala 30:26]
  wire [607:0] meta_s_axis_tdata; // @[Meta.scala 30:26]
  wire  meta_s_axis_tdest; // @[Meta.scala 30:26]
  wire  meta_s_axis_tid; // @[Meta.scala 30:26]
  wire [75:0] meta_s_axis_tkeep; // @[Meta.scala 30:26]
  wire  meta_s_axis_tlast; // @[Meta.scala 30:26]
  wire [75:0] meta_s_axis_tstrb; // @[Meta.scala 30:26]
  wire  meta_s_axis_tuser; // @[Meta.scala 30:26]
  wire  meta_s_axis_tvalid; // @[Meta.scala 30:26]
  xpm_fifo_axis
    #(.RD_DATA_COUNT_WIDTH(5), .CLOCKING_MODE("independent_clock"), .PACKET_FIFO("false"), .USE_ADV_FEATURES("0404"), .TID_WIDTH(1), .TDEST_WIDTH(1), .PROG_EMPTY_THRESH(10), .TUSER_WIDTH(1), .FIFO_DEPTH(16), .SIM_ASSERT_CHK(0), .WR_DATA_COUNT_WIDTH(5), .ECC_MODE("no_ecc"), .FIFO_MEMORY_TYPE("auto"), .PROG_FULL_THRESH(10), .TDATA_WIDTH(608), .RELATED_CLOCKS(0), .CASCADE_HEIGHT(0), .CDC_SYNC_STAGES(2))
    meta ( // @[Meta.scala 30:26]
    .m_axis_tdata(meta_m_axis_tdata),
    .m_axis_tkeep(meta_m_axis_tkeep),
    .m_axis_tlast(meta_m_axis_tlast),
    .m_axis_tvalid(meta_m_axis_tvalid),
    .rd_data_count_axis(meta_rd_data_count_axis),
    .s_axis_tready(meta_s_axis_tready),
    .wr_data_count_axis(meta_wr_data_count_axis),
    .m_aclk(meta_m_aclk),
    .m_axis_tready(meta_m_axis_tready),
    .s_aclk(meta_s_aclk),
    .s_aresetn(meta_s_aresetn),
    .s_axis_tdata(meta_s_axis_tdata),
    .s_axis_tdest(meta_s_axis_tdest),
    .s_axis_tid(meta_s_axis_tid),
    .s_axis_tkeep(meta_s_axis_tkeep),
    .s_axis_tlast(meta_s_axis_tlast),
    .s_axis_tstrb(meta_s_axis_tstrb),
    .s_axis_tuser(meta_s_axis_tuser),
    .s_axis_tvalid(meta_s_axis_tvalid)
  );
  assign io_in_ready = meta_s_axis_tready; // @[Meta.scala 34:41]
  assign io_out_data = meta_m_axis_tdata; // @[Meta.scala 31:41]
  assign io_out_valid = meta_m_axis_tvalid; // @[Meta.scala 32:41]
  assign meta_m_aclk = io_m_clk; // @[Meta.scala 37:49]
  assign meta_m_axis_tready = io_out_ready; // @[Meta.scala 38:41]
  assign meta_s_aclk = io_s_clk; // @[Meta.scala 39:49]
  assign meta_s_aresetn = io_reset_n; // @[Meta.scala 40:49]
  assign meta_s_axis_tdata = io_in_data; // @[Meta.scala 41:41]
  assign meta_s_axis_tdest = 1'h0; // @[Meta.scala 42:41]
  assign meta_s_axis_tid = 1'h0; // @[Meta.scala 43:49]
  assign meta_s_axis_tkeep = 76'hfffffffffffffffffff; // @[Bitwise.scala 72:12]
  assign meta_s_axis_tlast = 1'h1; // @[Meta.scala 45:41]
  assign meta_s_axis_tstrb = 76'hfffffffffffffffffff; // @[Bitwise.scala 72:12]
  assign meta_s_axis_tuser = 1'h0; // @[Meta.scala 47:41]
  assign meta_s_axis_tvalid = io_in_valid; // @[Meta.scala 48:41]
endmodule
module XConverter_1(
  input          io__in_clk,
  input          io__out_clk,
  input          io__rstn,
  output         io__in_ready,
  input          io__in_valid,
  input  [511:0] io__in_bits_data,
  input  [31:0]  io__in_bits_tcrc,
  input          io__in_bits_ctrl_marker,
  input  [6:0]   io__in_bits_ctrl_ecc,
  input  [31:0]  io__in_bits_ctrl_len,
  input  [2:0]   io__in_bits_ctrl_port_id,
  input  [10:0]  io__in_bits_ctrl_qid,
  input          io__in_bits_ctrl_has_cmpt,
  input          io__in_bits_last,
  input  [5:0]   io__in_bits_mty,
  input          io__out_ready,
  output         io__out_valid,
  output [511:0] io__out_bits_data,
  output [31:0]  io__out_bits_tcrc,
  output         io__out_bits_ctrl_marker,
  output [6:0]   io__out_bits_ctrl_ecc,
  output [31:0]  io__out_bits_ctrl_len,
  output [2:0]   io__out_bits_ctrl_port_id,
  output [10:0]  io__out_bits_ctrl_qid,
  output         io__out_bits_ctrl_has_cmpt,
  output         io__out_bits_last,
  output [5:0]   io__out_bits_mty,
  output         io_out_ready,
  output         io_out_valid_0
);
  wire  fifo_io_m_clk; // @[XConverter.scala 97:34]
  wire  fifo_io_s_clk; // @[XConverter.scala 97:34]
  wire  fifo_io_reset_n; // @[XConverter.scala 97:34]
  wire [607:0] fifo_io_in_data; // @[XConverter.scala 97:34]
  wire  fifo_io_in_valid; // @[XConverter.scala 97:34]
  wire  fifo_io_in_ready; // @[XConverter.scala 97:34]
  wire [607:0] fifo_io_out_data; // @[XConverter.scala 97:34]
  wire  fifo_io_out_valid; // @[XConverter.scala 97:34]
  wire  fifo_io_out_ready; // @[XConverter.scala 97:34]
  wire [605:0] _fifo_io_in_data_T = {io__in_bits_data,io__in_bits_tcrc,io__in_bits_ctrl_marker,io__in_bits_ctrl_ecc,
    io__in_bits_ctrl_len,io__in_bits_ctrl_port_id,io__in_bits_ctrl_qid,io__in_bits_ctrl_has_cmpt,io__in_bits_last,
    io__in_bits_mty}; // @[XConverter.scala 103:63]
  SV_STREAM_FIFO_1 fifo ( // @[XConverter.scala 97:34]
    .io_m_clk(fifo_io_m_clk),
    .io_s_clk(fifo_io_s_clk),
    .io_reset_n(fifo_io_reset_n),
    .io_in_data(fifo_io_in_data),
    .io_in_valid(fifo_io_in_valid),
    .io_in_ready(fifo_io_in_ready),
    .io_out_data(fifo_io_out_data),
    .io_out_valid(fifo_io_out_valid),
    .io_out_ready(fifo_io_out_ready)
  );
  assign io__in_ready = fifo_io_in_ready; // @[XConverter.scala 105:41]
  assign io__out_valid = fifo_io_out_valid; // @[XConverter.scala 108:41]
  assign io__out_bits_data = fifo_io_out_data[605:94]; // @[XConverter.scala 107:77]
  assign io__out_bits_tcrc = fifo_io_out_data[93:62]; // @[XConverter.scala 107:77]
  assign io__out_bits_ctrl_marker = fifo_io_out_data[61]; // @[XConverter.scala 107:77]
  assign io__out_bits_ctrl_ecc = fifo_io_out_data[60:54]; // @[XConverter.scala 107:77]
  assign io__out_bits_ctrl_len = fifo_io_out_data[53:22]; // @[XConverter.scala 107:77]
  assign io__out_bits_ctrl_port_id = fifo_io_out_data[21:19]; // @[XConverter.scala 107:77]
  assign io__out_bits_ctrl_qid = fifo_io_out_data[18:8]; // @[XConverter.scala 107:77]
  assign io__out_bits_ctrl_has_cmpt = fifo_io_out_data[7]; // @[XConverter.scala 107:77]
  assign io__out_bits_last = fifo_io_out_data[6]; // @[XConverter.scala 107:77]
  assign io__out_bits_mty = fifo_io_out_data[5:0]; // @[XConverter.scala 107:77]
  assign io_out_ready = io__out_ready;
  assign io_out_valid_0 = io__out_valid;
  assign fifo_io_m_clk = io__out_clk; // @[XConverter.scala 100:41]
  assign fifo_io_s_clk = io__in_clk; // @[XConverter.scala 99:41]
  assign fifo_io_reset_n = io__rstn; // @[XConverter.scala 101:41]
  assign fifo_io_in_data = {{2'd0}, _fifo_io_in_data_T}; // @[XConverter.scala 103:63]
  assign fifo_io_in_valid = io__in_valid; // @[XConverter.scala 104:41]
  assign fifo_io_out_ready = io__out_ready; // @[XConverter.scala 109:41]
endmodule
module RegSlice_1(
  input          clock,
  input          reset,
  output         io_upStream_ready,
  input          io_upStream_valid,
  input  [511:0] io_upStream_bits_data,
  input  [31:0]  io_upStream_bits_tcrc,
  input          io_upStream_bits_ctrl_marker,
  input  [6:0]   io_upStream_bits_ctrl_ecc,
  input  [31:0]  io_upStream_bits_ctrl_len,
  input  [2:0]   io_upStream_bits_ctrl_port_id,
  input  [10:0]  io_upStream_bits_ctrl_qid,
  input          io_upStream_bits_ctrl_has_cmpt,
  input          io_upStream_bits_last,
  input  [5:0]   io_upStream_bits_mty,
  input          io_downStream_ready,
  output         io_downStream_valid,
  output [511:0] io_downStream_bits_data,
  output [31:0]  io_downStream_bits_tcrc,
  output         io_downStream_bits_ctrl_marker,
  output [6:0]   io_downStream_bits_ctrl_ecc,
  output [31:0]  io_downStream_bits_ctrl_len,
  output [2:0]   io_downStream_bits_ctrl_port_id,
  output [10:0]  io_downStream_bits_ctrl_qid,
  output         io_downStream_bits_ctrl_has_cmpt,
  output         io_downStream_bits_last,
  output [5:0]   io_downStream_bits_mty
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [511:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [511:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
`endif // RANDOMIZE_REG_INIT
  reg  fwd_valid; // @[RegSlices.scala 112:34]
  reg [511:0] fwd_data_data; // @[RegSlices.scala 113:30]
  reg [31:0] fwd_data_tcrc; // @[RegSlices.scala 113:30]
  reg  fwd_data_ctrl_marker; // @[RegSlices.scala 113:30]
  reg [6:0] fwd_data_ctrl_ecc; // @[RegSlices.scala 113:30]
  reg [31:0] fwd_data_ctrl_len; // @[RegSlices.scala 113:30]
  reg [2:0] fwd_data_ctrl_port_id; // @[RegSlices.scala 113:30]
  reg [10:0] fwd_data_ctrl_qid; // @[RegSlices.scala 113:30]
  reg  fwd_data_ctrl_has_cmpt; // @[RegSlices.scala 113:30]
  reg  fwd_data_last; // @[RegSlices.scala 113:30]
  reg [5:0] fwd_data_mty; // @[RegSlices.scala 113:30]
  wire  fwd_ready_s = ~fwd_valid | io_downStream_ready; // @[RegSlices.scala 115:35]
  reg  bwd_ready; // @[RegSlices.scala 123:34]
  reg [511:0] bwd_data_data; // @[RegSlices.scala 124:30]
  reg [31:0] bwd_data_tcrc; // @[RegSlices.scala 124:30]
  reg  bwd_data_ctrl_marker; // @[RegSlices.scala 124:30]
  reg [6:0] bwd_data_ctrl_ecc; // @[RegSlices.scala 124:30]
  reg [31:0] bwd_data_ctrl_len; // @[RegSlices.scala 124:30]
  reg [2:0] bwd_data_ctrl_port_id; // @[RegSlices.scala 124:30]
  reg [10:0] bwd_data_ctrl_qid; // @[RegSlices.scala 124:30]
  reg  bwd_data_ctrl_has_cmpt; // @[RegSlices.scala 124:30]
  reg  bwd_data_last; // @[RegSlices.scala 124:30]
  reg [5:0] bwd_data_mty; // @[RegSlices.scala 124:30]
  wire  _fwd_valid_T = io_downStream_ready ? 1'h0 : fwd_valid; // @[RegSlices.scala 121:53]
  wire  bwd_valid_s = ~bwd_ready | io_upStream_valid; // @[RegSlices.scala 126:39]
  wire  _bwd_ready_T = io_upStream_valid ? 1'h0 : bwd_ready; // @[RegSlices.scala 132:53]
  assign io_upStream_ready = bwd_ready; // @[RegSlices.scala 107:31 RegSlices.scala 128:25]
  assign io_downStream_valid = fwd_valid; // @[RegSlices.scala 109:31 RegSlices.scala 116:21]
  assign io_downStream_bits_data = fwd_data_data; // @[RegSlices.scala 108:31 RegSlices.scala 117:25]
  assign io_downStream_bits_tcrc = fwd_data_tcrc; // @[RegSlices.scala 108:31 RegSlices.scala 117:25]
  assign io_downStream_bits_ctrl_marker = fwd_data_ctrl_marker; // @[RegSlices.scala 108:31 RegSlices.scala 117:25]
  assign io_downStream_bits_ctrl_ecc = fwd_data_ctrl_ecc; // @[RegSlices.scala 108:31 RegSlices.scala 117:25]
  assign io_downStream_bits_ctrl_len = fwd_data_ctrl_len; // @[RegSlices.scala 108:31 RegSlices.scala 117:25]
  assign io_downStream_bits_ctrl_port_id = fwd_data_ctrl_port_id; // @[RegSlices.scala 108:31 RegSlices.scala 117:25]
  assign io_downStream_bits_ctrl_qid = fwd_data_ctrl_qid; // @[RegSlices.scala 108:31 RegSlices.scala 117:25]
  assign io_downStream_bits_ctrl_has_cmpt = fwd_data_ctrl_has_cmpt; // @[RegSlices.scala 108:31 RegSlices.scala 117:25]
  assign io_downStream_bits_last = fwd_data_last; // @[RegSlices.scala 108:31 RegSlices.scala 117:25]
  assign io_downStream_bits_mty = fwd_data_mty; // @[RegSlices.scala 108:31 RegSlices.scala 117:25]
  always @(posedge clock) begin
    if (reset) begin // @[RegSlices.scala 112:34]
      fwd_valid <= 1'h0; // @[RegSlices.scala 112:34]
    end else begin
      fwd_valid <= bwd_valid_s | _fwd_valid_T; // @[RegSlices.scala 121:25]
    end
    if (fwd_ready_s) begin // @[RegSlices.scala 119:31]
      if (bwd_ready) begin // @[RegSlices.scala 127:31]
        fwd_data_data <= io_upStream_bits_data;
      end else begin
        fwd_data_data <= bwd_data_data;
      end
    end
    if (fwd_ready_s) begin // @[RegSlices.scala 119:31]
      if (bwd_ready) begin // @[RegSlices.scala 127:31]
        fwd_data_tcrc <= io_upStream_bits_tcrc;
      end else begin
        fwd_data_tcrc <= bwd_data_tcrc;
      end
    end
    if (fwd_ready_s) begin // @[RegSlices.scala 119:31]
      if (bwd_ready) begin // @[RegSlices.scala 127:31]
        fwd_data_ctrl_marker <= io_upStream_bits_ctrl_marker;
      end else begin
        fwd_data_ctrl_marker <= bwd_data_ctrl_marker;
      end
    end
    if (fwd_ready_s) begin // @[RegSlices.scala 119:31]
      if (bwd_ready) begin // @[RegSlices.scala 127:31]
        fwd_data_ctrl_ecc <= io_upStream_bits_ctrl_ecc;
      end else begin
        fwd_data_ctrl_ecc <= bwd_data_ctrl_ecc;
      end
    end
    if (fwd_ready_s) begin // @[RegSlices.scala 119:31]
      if (bwd_ready) begin // @[RegSlices.scala 127:31]
        fwd_data_ctrl_len <= io_upStream_bits_ctrl_len;
      end else begin
        fwd_data_ctrl_len <= bwd_data_ctrl_len;
      end
    end
    if (fwd_ready_s) begin // @[RegSlices.scala 119:31]
      if (bwd_ready) begin // @[RegSlices.scala 127:31]
        fwd_data_ctrl_port_id <= io_upStream_bits_ctrl_port_id;
      end else begin
        fwd_data_ctrl_port_id <= bwd_data_ctrl_port_id;
      end
    end
    if (fwd_ready_s) begin // @[RegSlices.scala 119:31]
      if (bwd_ready) begin // @[RegSlices.scala 127:31]
        fwd_data_ctrl_qid <= io_upStream_bits_ctrl_qid;
      end else begin
        fwd_data_ctrl_qid <= bwd_data_ctrl_qid;
      end
    end
    if (fwd_ready_s) begin // @[RegSlices.scala 119:31]
      if (bwd_ready) begin // @[RegSlices.scala 127:31]
        fwd_data_ctrl_has_cmpt <= io_upStream_bits_ctrl_has_cmpt;
      end else begin
        fwd_data_ctrl_has_cmpt <= bwd_data_ctrl_has_cmpt;
      end
    end
    if (fwd_ready_s) begin // @[RegSlices.scala 119:31]
      if (bwd_ready) begin // @[RegSlices.scala 127:31]
        fwd_data_last <= io_upStream_bits_last;
      end else begin
        fwd_data_last <= bwd_data_last;
      end
    end
    if (fwd_ready_s) begin // @[RegSlices.scala 119:31]
      if (bwd_ready) begin // @[RegSlices.scala 127:31]
        fwd_data_mty <= io_upStream_bits_mty;
      end else begin
        fwd_data_mty <= bwd_data_mty;
      end
    end
    bwd_ready <= reset | (fwd_ready_s | _bwd_ready_T); // @[RegSlices.scala 123:34 RegSlices.scala 123:34 RegSlices.scala 132:25]
    if (bwd_ready) begin // @[RegSlices.scala 130:31]
      bwd_data_data <= io_upStream_bits_data;
    end
    if (bwd_ready) begin // @[RegSlices.scala 130:31]
      bwd_data_tcrc <= io_upStream_bits_tcrc;
    end
    if (bwd_ready) begin // @[RegSlices.scala 130:31]
      bwd_data_ctrl_marker <= io_upStream_bits_ctrl_marker;
    end
    if (bwd_ready) begin // @[RegSlices.scala 130:31]
      bwd_data_ctrl_ecc <= io_upStream_bits_ctrl_ecc;
    end
    if (bwd_ready) begin // @[RegSlices.scala 130:31]
      bwd_data_ctrl_len <= io_upStream_bits_ctrl_len;
    end
    if (bwd_ready) begin // @[RegSlices.scala 130:31]
      bwd_data_ctrl_port_id <= io_upStream_bits_ctrl_port_id;
    end
    if (bwd_ready) begin // @[RegSlices.scala 130:31]
      bwd_data_ctrl_qid <= io_upStream_bits_ctrl_qid;
    end
    if (bwd_ready) begin // @[RegSlices.scala 130:31]
      bwd_data_ctrl_has_cmpt <= io_upStream_bits_ctrl_has_cmpt;
    end
    if (bwd_ready) begin // @[RegSlices.scala 130:31]
      bwd_data_last <= io_upStream_bits_last;
    end
    if (bwd_ready) begin // @[RegSlices.scala 130:31]
      bwd_data_mty <= io_upStream_bits_mty;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  fwd_valid = _RAND_0[0:0];
  _RAND_1 = {16{`RANDOM}};
  fwd_data_data = _RAND_1[511:0];
  _RAND_2 = {1{`RANDOM}};
  fwd_data_tcrc = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  fwd_data_ctrl_marker = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  fwd_data_ctrl_ecc = _RAND_4[6:0];
  _RAND_5 = {1{`RANDOM}};
  fwd_data_ctrl_len = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  fwd_data_ctrl_port_id = _RAND_6[2:0];
  _RAND_7 = {1{`RANDOM}};
  fwd_data_ctrl_qid = _RAND_7[10:0];
  _RAND_8 = {1{`RANDOM}};
  fwd_data_ctrl_has_cmpt = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  fwd_data_last = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  fwd_data_mty = _RAND_10[5:0];
  _RAND_11 = {1{`RANDOM}};
  bwd_ready = _RAND_11[0:0];
  _RAND_12 = {16{`RANDOM}};
  bwd_data_data = _RAND_12[511:0];
  _RAND_13 = {1{`RANDOM}};
  bwd_data_tcrc = _RAND_13[31:0];
  _RAND_14 = {1{`RANDOM}};
  bwd_data_ctrl_marker = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  bwd_data_ctrl_ecc = _RAND_15[6:0];
  _RAND_16 = {1{`RANDOM}};
  bwd_data_ctrl_len = _RAND_16[31:0];
  _RAND_17 = {1{`RANDOM}};
  bwd_data_ctrl_port_id = _RAND_17[2:0];
  _RAND_18 = {1{`RANDOM}};
  bwd_data_ctrl_qid = _RAND_18[10:0];
  _RAND_19 = {1{`RANDOM}};
  bwd_data_ctrl_has_cmpt = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  bwd_data_last = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  bwd_data_mty = _RAND_21[5:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module SV_STREAM_FIFO_2(
  input          io_m_clk,
  input          io_s_clk,
  input          io_reset_n,
  input  [143:0] io_in_data,
  input          io_in_valid,
  output         io_in_ready,
  output [143:0] io_out_data,
  output         io_out_valid,
  input          io_out_ready
);
  wire [143:0] meta_m_axis_tdata; // @[Meta.scala 30:26]
  wire [17:0] meta_m_axis_tkeep; // @[Meta.scala 30:26]
  wire  meta_m_axis_tlast; // @[Meta.scala 30:26]
  wire  meta_m_axis_tvalid; // @[Meta.scala 30:26]
  wire [4:0] meta_rd_data_count_axis; // @[Meta.scala 30:26]
  wire  meta_s_axis_tready; // @[Meta.scala 30:26]
  wire [4:0] meta_wr_data_count_axis; // @[Meta.scala 30:26]
  wire  meta_m_aclk; // @[Meta.scala 30:26]
  wire  meta_m_axis_tready; // @[Meta.scala 30:26]
  wire  meta_s_aclk; // @[Meta.scala 30:26]
  wire  meta_s_aresetn; // @[Meta.scala 30:26]
  wire [143:0] meta_s_axis_tdata; // @[Meta.scala 30:26]
  wire  meta_s_axis_tdest; // @[Meta.scala 30:26]
  wire  meta_s_axis_tid; // @[Meta.scala 30:26]
  wire [17:0] meta_s_axis_tkeep; // @[Meta.scala 30:26]
  wire  meta_s_axis_tlast; // @[Meta.scala 30:26]
  wire [17:0] meta_s_axis_tstrb; // @[Meta.scala 30:26]
  wire  meta_s_axis_tuser; // @[Meta.scala 30:26]
  wire  meta_s_axis_tvalid; // @[Meta.scala 30:26]
  xpm_fifo_axis
    #(.RD_DATA_COUNT_WIDTH(5), .CLOCKING_MODE("independent_clock"), .PACKET_FIFO("false"), .USE_ADV_FEATURES("0404"), .TID_WIDTH(1), .TDEST_WIDTH(1), .PROG_EMPTY_THRESH(10), .TUSER_WIDTH(1), .FIFO_DEPTH(16), .SIM_ASSERT_CHK(0), .WR_DATA_COUNT_WIDTH(5), .ECC_MODE("no_ecc"), .FIFO_MEMORY_TYPE("auto"), .PROG_FULL_THRESH(10), .TDATA_WIDTH(144), .RELATED_CLOCKS(0), .CASCADE_HEIGHT(0), .CDC_SYNC_STAGES(2))
    meta ( // @[Meta.scala 30:26]
    .m_axis_tdata(meta_m_axis_tdata),
    .m_axis_tkeep(meta_m_axis_tkeep),
    .m_axis_tlast(meta_m_axis_tlast),
    .m_axis_tvalid(meta_m_axis_tvalid),
    .rd_data_count_axis(meta_rd_data_count_axis),
    .s_axis_tready(meta_s_axis_tready),
    .wr_data_count_axis(meta_wr_data_count_axis),
    .m_aclk(meta_m_aclk),
    .m_axis_tready(meta_m_axis_tready),
    .s_aclk(meta_s_aclk),
    .s_aresetn(meta_s_aresetn),
    .s_axis_tdata(meta_s_axis_tdata),
    .s_axis_tdest(meta_s_axis_tdest),
    .s_axis_tid(meta_s_axis_tid),
    .s_axis_tkeep(meta_s_axis_tkeep),
    .s_axis_tlast(meta_s_axis_tlast),
    .s_axis_tstrb(meta_s_axis_tstrb),
    .s_axis_tuser(meta_s_axis_tuser),
    .s_axis_tvalid(meta_s_axis_tvalid)
  );
  assign io_in_ready = meta_s_axis_tready; // @[Meta.scala 34:41]
  assign io_out_data = meta_m_axis_tdata; // @[Meta.scala 31:41]
  assign io_out_valid = meta_m_axis_tvalid; // @[Meta.scala 32:41]
  assign meta_m_aclk = io_m_clk; // @[Meta.scala 37:49]
  assign meta_m_axis_tready = io_out_ready; // @[Meta.scala 38:41]
  assign meta_s_aclk = io_s_clk; // @[Meta.scala 39:49]
  assign meta_s_aresetn = io_reset_n; // @[Meta.scala 40:49]
  assign meta_s_axis_tdata = io_in_data; // @[Meta.scala 41:41]
  assign meta_s_axis_tdest = 1'h0; // @[Meta.scala 42:41]
  assign meta_s_axis_tid = 1'h0; // @[Meta.scala 43:49]
  assign meta_s_axis_tkeep = 18'h3ffff; // @[Bitwise.scala 72:12]
  assign meta_s_axis_tlast = 1'h1; // @[Meta.scala 45:41]
  assign meta_s_axis_tstrb = 18'h3ffff; // @[Bitwise.scala 72:12]
  assign meta_s_axis_tuser = 1'h0; // @[Meta.scala 47:41]
  assign meta_s_axis_tvalid = io_in_valid; // @[Meta.scala 48:41]
endmodule
module XConverter_2(
  input         io__in_clk,
  input         io__out_clk,
  input         io__rstn,
  output        io__in_ready,
  input         io__in_valid,
  input  [63:0] io__in_bits_addr,
  input  [31:0] io__in_bits_len,
  input         io__in_bits_eop,
  input         io__in_bits_sop,
  input         io__in_bits_mrkr_req,
  input         io__in_bits_sdi,
  input  [10:0] io__in_bits_qid,
  input         io__in_bits_error,
  input  [7:0]  io__in_bits_func,
  input  [15:0] io__in_bits_cidx,
  input  [2:0]  io__in_bits_port_id,
  input         io__in_bits_no_dma,
  input         io__out_ready,
  output        io__out_valid,
  output [63:0] io__out_bits_addr,
  output [31:0] io__out_bits_len,
  output        io__out_bits_eop,
  output        io__out_bits_sop,
  output        io__out_bits_mrkr_req,
  output        io__out_bits_sdi,
  output [10:0] io__out_bits_qid,
  output        io__out_bits_error,
  output [7:0]  io__out_bits_func,
  output [15:0] io__out_bits_cidx,
  output [2:0]  io__out_bits_port_id,
  output        io__out_bits_no_dma,
  output        io_out_valid,
  output        io_out_ready_1
);
  wire  fifo_io_m_clk; // @[XConverter.scala 97:34]
  wire  fifo_io_s_clk; // @[XConverter.scala 97:34]
  wire  fifo_io_reset_n; // @[XConverter.scala 97:34]
  wire [143:0] fifo_io_in_data; // @[XConverter.scala 97:34]
  wire  fifo_io_in_valid; // @[XConverter.scala 97:34]
  wire  fifo_io_in_ready; // @[XConverter.scala 97:34]
  wire [143:0] fifo_io_out_data; // @[XConverter.scala 97:34]
  wire  fifo_io_out_valid; // @[XConverter.scala 97:34]
  wire  fifo_io_out_ready; // @[XConverter.scala 97:34]
  wire [39:0] fifo_io_in_data_lo = {io__in_bits_qid,io__in_bits_error,io__in_bits_func,io__in_bits_cidx,
    io__in_bits_port_id,io__in_bits_no_dma}; // @[XConverter.scala 103:63]
  wire [139:0] _fifo_io_in_data_T = {io__in_bits_addr,io__in_bits_len,io__in_bits_eop,io__in_bits_sop,
    io__in_bits_mrkr_req,io__in_bits_sdi,fifo_io_in_data_lo}; // @[XConverter.scala 103:63]
  SV_STREAM_FIFO_2 fifo ( // @[XConverter.scala 97:34]
    .io_m_clk(fifo_io_m_clk),
    .io_s_clk(fifo_io_s_clk),
    .io_reset_n(fifo_io_reset_n),
    .io_in_data(fifo_io_in_data),
    .io_in_valid(fifo_io_in_valid),
    .io_in_ready(fifo_io_in_ready),
    .io_out_data(fifo_io_out_data),
    .io_out_valid(fifo_io_out_valid),
    .io_out_ready(fifo_io_out_ready)
  );
  assign io__in_ready = fifo_io_in_ready; // @[XConverter.scala 105:41]
  assign io__out_valid = fifo_io_out_valid; // @[XConverter.scala 108:41]
  assign io__out_bits_addr = fifo_io_out_data[139:76]; // @[XConverter.scala 107:77]
  assign io__out_bits_len = fifo_io_out_data[75:44]; // @[XConverter.scala 107:77]
  assign io__out_bits_eop = fifo_io_out_data[43]; // @[XConverter.scala 107:77]
  assign io__out_bits_sop = fifo_io_out_data[42]; // @[XConverter.scala 107:77]
  assign io__out_bits_mrkr_req = fifo_io_out_data[41]; // @[XConverter.scala 107:77]
  assign io__out_bits_sdi = fifo_io_out_data[40]; // @[XConverter.scala 107:77]
  assign io__out_bits_qid = fifo_io_out_data[39:29]; // @[XConverter.scala 107:77]
  assign io__out_bits_error = fifo_io_out_data[28]; // @[XConverter.scala 107:77]
  assign io__out_bits_func = fifo_io_out_data[27:20]; // @[XConverter.scala 107:77]
  assign io__out_bits_cidx = fifo_io_out_data[19:4]; // @[XConverter.scala 107:77]
  assign io__out_bits_port_id = fifo_io_out_data[3:1]; // @[XConverter.scala 107:77]
  assign io__out_bits_no_dma = fifo_io_out_data[0]; // @[XConverter.scala 107:77]
  assign io_out_valid = io__out_valid;
  assign io_out_ready_1 = io__out_ready;
  assign fifo_io_m_clk = io__out_clk; // @[XConverter.scala 100:41]
  assign fifo_io_s_clk = io__in_clk; // @[XConverter.scala 99:41]
  assign fifo_io_reset_n = io__rstn; // @[XConverter.scala 101:41]
  assign fifo_io_in_data = {{4'd0}, _fifo_io_in_data_T}; // @[XConverter.scala 103:63]
  assign fifo_io_in_valid = io__in_valid; // @[XConverter.scala 104:41]
  assign fifo_io_out_ready = io__out_ready; // @[XConverter.scala 109:41]
endmodule
module RegSlice_2(
  input         clock,
  input         reset,
  output        io_upStream_ready,
  input         io_upStream_valid,
  input  [63:0] io_upStream_bits_addr,
  input  [31:0] io_upStream_bits_len,
  input         io_upStream_bits_eop,
  input         io_upStream_bits_sop,
  input         io_upStream_bits_mrkr_req,
  input         io_upStream_bits_sdi,
  input  [10:0] io_upStream_bits_qid,
  input         io_upStream_bits_error,
  input  [7:0]  io_upStream_bits_func,
  input  [15:0] io_upStream_bits_cidx,
  input  [2:0]  io_upStream_bits_port_id,
  input         io_upStream_bits_no_dma,
  input         io_downStream_ready,
  output        io_downStream_valid,
  output [63:0] io_downStream_bits_addr,
  output [31:0] io_downStream_bits_len,
  output        io_downStream_bits_eop,
  output        io_downStream_bits_sop,
  output        io_downStream_bits_mrkr_req,
  output        io_downStream_bits_sdi,
  output [10:0] io_downStream_bits_qid,
  output        io_downStream_bits_error,
  output [7:0]  io_downStream_bits_func,
  output [15:0] io_downStream_bits_cidx,
  output [2:0]  io_downStream_bits_port_id,
  output        io_downStream_bits_no_dma
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [63:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
`endif // RANDOMIZE_REG_INIT
  reg  fwd_valid; // @[RegSlices.scala 112:34]
  reg [63:0] fwd_data_addr; // @[RegSlices.scala 113:30]
  reg [31:0] fwd_data_len; // @[RegSlices.scala 113:30]
  reg  fwd_data_eop; // @[RegSlices.scala 113:30]
  reg  fwd_data_sop; // @[RegSlices.scala 113:30]
  reg  fwd_data_mrkr_req; // @[RegSlices.scala 113:30]
  reg  fwd_data_sdi; // @[RegSlices.scala 113:30]
  reg [10:0] fwd_data_qid; // @[RegSlices.scala 113:30]
  reg  fwd_data_error; // @[RegSlices.scala 113:30]
  reg [7:0] fwd_data_func; // @[RegSlices.scala 113:30]
  reg [15:0] fwd_data_cidx; // @[RegSlices.scala 113:30]
  reg [2:0] fwd_data_port_id; // @[RegSlices.scala 113:30]
  reg  fwd_data_no_dma; // @[RegSlices.scala 113:30]
  wire  fwd_ready_s = ~fwd_valid | io_downStream_ready; // @[RegSlices.scala 115:35]
  reg  bwd_ready; // @[RegSlices.scala 123:34]
  reg [63:0] bwd_data_addr; // @[RegSlices.scala 124:30]
  reg [31:0] bwd_data_len; // @[RegSlices.scala 124:30]
  reg  bwd_data_eop; // @[RegSlices.scala 124:30]
  reg  bwd_data_sop; // @[RegSlices.scala 124:30]
  reg  bwd_data_mrkr_req; // @[RegSlices.scala 124:30]
  reg  bwd_data_sdi; // @[RegSlices.scala 124:30]
  reg [10:0] bwd_data_qid; // @[RegSlices.scala 124:30]
  reg  bwd_data_error; // @[RegSlices.scala 124:30]
  reg [7:0] bwd_data_func; // @[RegSlices.scala 124:30]
  reg [15:0] bwd_data_cidx; // @[RegSlices.scala 124:30]
  reg [2:0] bwd_data_port_id; // @[RegSlices.scala 124:30]
  reg  bwd_data_no_dma; // @[RegSlices.scala 124:30]
  wire  _fwd_valid_T = io_downStream_ready ? 1'h0 : fwd_valid; // @[RegSlices.scala 121:53]
  wire  bwd_valid_s = ~bwd_ready | io_upStream_valid; // @[RegSlices.scala 126:39]
  wire  _bwd_ready_T = io_upStream_valid ? 1'h0 : bwd_ready; // @[RegSlices.scala 132:53]
  assign io_upStream_ready = bwd_ready; // @[RegSlices.scala 107:31 RegSlices.scala 128:25]
  assign io_downStream_valid = fwd_valid; // @[RegSlices.scala 109:31 RegSlices.scala 116:21]
  assign io_downStream_bits_addr = fwd_data_addr; // @[RegSlices.scala 108:31 RegSlices.scala 117:25]
  assign io_downStream_bits_len = fwd_data_len; // @[RegSlices.scala 108:31 RegSlices.scala 117:25]
  assign io_downStream_bits_eop = fwd_data_eop; // @[RegSlices.scala 108:31 RegSlices.scala 117:25]
  assign io_downStream_bits_sop = fwd_data_sop; // @[RegSlices.scala 108:31 RegSlices.scala 117:25]
  assign io_downStream_bits_mrkr_req = fwd_data_mrkr_req; // @[RegSlices.scala 108:31 RegSlices.scala 117:25]
  assign io_downStream_bits_sdi = fwd_data_sdi; // @[RegSlices.scala 108:31 RegSlices.scala 117:25]
  assign io_downStream_bits_qid = fwd_data_qid; // @[RegSlices.scala 108:31 RegSlices.scala 117:25]
  assign io_downStream_bits_error = fwd_data_error; // @[RegSlices.scala 108:31 RegSlices.scala 117:25]
  assign io_downStream_bits_func = fwd_data_func; // @[RegSlices.scala 108:31 RegSlices.scala 117:25]
  assign io_downStream_bits_cidx = fwd_data_cidx; // @[RegSlices.scala 108:31 RegSlices.scala 117:25]
  assign io_downStream_bits_port_id = fwd_data_port_id; // @[RegSlices.scala 108:31 RegSlices.scala 117:25]
  assign io_downStream_bits_no_dma = fwd_data_no_dma; // @[RegSlices.scala 108:31 RegSlices.scala 117:25]
  always @(posedge clock) begin
    if (reset) begin // @[RegSlices.scala 112:34]
      fwd_valid <= 1'h0; // @[RegSlices.scala 112:34]
    end else begin
      fwd_valid <= bwd_valid_s | _fwd_valid_T; // @[RegSlices.scala 121:25]
    end
    if (fwd_ready_s) begin // @[RegSlices.scala 119:31]
      if (bwd_ready) begin // @[RegSlices.scala 127:31]
        fwd_data_addr <= io_upStream_bits_addr;
      end else begin
        fwd_data_addr <= bwd_data_addr;
      end
    end
    if (fwd_ready_s) begin // @[RegSlices.scala 119:31]
      if (bwd_ready) begin // @[RegSlices.scala 127:31]
        fwd_data_len <= io_upStream_bits_len;
      end else begin
        fwd_data_len <= bwd_data_len;
      end
    end
    if (fwd_ready_s) begin // @[RegSlices.scala 119:31]
      if (bwd_ready) begin // @[RegSlices.scala 127:31]
        fwd_data_eop <= io_upStream_bits_eop;
      end else begin
        fwd_data_eop <= bwd_data_eop;
      end
    end
    if (fwd_ready_s) begin // @[RegSlices.scala 119:31]
      if (bwd_ready) begin // @[RegSlices.scala 127:31]
        fwd_data_sop <= io_upStream_bits_sop;
      end else begin
        fwd_data_sop <= bwd_data_sop;
      end
    end
    if (fwd_ready_s) begin // @[RegSlices.scala 119:31]
      if (bwd_ready) begin // @[RegSlices.scala 127:31]
        fwd_data_mrkr_req <= io_upStream_bits_mrkr_req;
      end else begin
        fwd_data_mrkr_req <= bwd_data_mrkr_req;
      end
    end
    if (fwd_ready_s) begin // @[RegSlices.scala 119:31]
      if (bwd_ready) begin // @[RegSlices.scala 127:31]
        fwd_data_sdi <= io_upStream_bits_sdi;
      end else begin
        fwd_data_sdi <= bwd_data_sdi;
      end
    end
    if (fwd_ready_s) begin // @[RegSlices.scala 119:31]
      if (bwd_ready) begin // @[RegSlices.scala 127:31]
        fwd_data_qid <= io_upStream_bits_qid;
      end else begin
        fwd_data_qid <= bwd_data_qid;
      end
    end
    if (fwd_ready_s) begin // @[RegSlices.scala 119:31]
      if (bwd_ready) begin // @[RegSlices.scala 127:31]
        fwd_data_error <= io_upStream_bits_error;
      end else begin
        fwd_data_error <= bwd_data_error;
      end
    end
    if (fwd_ready_s) begin // @[RegSlices.scala 119:31]
      if (bwd_ready) begin // @[RegSlices.scala 127:31]
        fwd_data_func <= io_upStream_bits_func;
      end else begin
        fwd_data_func <= bwd_data_func;
      end
    end
    if (fwd_ready_s) begin // @[RegSlices.scala 119:31]
      if (bwd_ready) begin // @[RegSlices.scala 127:31]
        fwd_data_cidx <= io_upStream_bits_cidx;
      end else begin
        fwd_data_cidx <= bwd_data_cidx;
      end
    end
    if (fwd_ready_s) begin // @[RegSlices.scala 119:31]
      if (bwd_ready) begin // @[RegSlices.scala 127:31]
        fwd_data_port_id <= io_upStream_bits_port_id;
      end else begin
        fwd_data_port_id <= bwd_data_port_id;
      end
    end
    if (fwd_ready_s) begin // @[RegSlices.scala 119:31]
      if (bwd_ready) begin // @[RegSlices.scala 127:31]
        fwd_data_no_dma <= io_upStream_bits_no_dma;
      end else begin
        fwd_data_no_dma <= bwd_data_no_dma;
      end
    end
    bwd_ready <= reset | (fwd_ready_s | _bwd_ready_T); // @[RegSlices.scala 123:34 RegSlices.scala 123:34 RegSlices.scala 132:25]
    if (bwd_ready) begin // @[RegSlices.scala 130:31]
      bwd_data_addr <= io_upStream_bits_addr;
    end
    if (bwd_ready) begin // @[RegSlices.scala 130:31]
      bwd_data_len <= io_upStream_bits_len;
    end
    if (bwd_ready) begin // @[RegSlices.scala 130:31]
      bwd_data_eop <= io_upStream_bits_eop;
    end
    if (bwd_ready) begin // @[RegSlices.scala 130:31]
      bwd_data_sop <= io_upStream_bits_sop;
    end
    if (bwd_ready) begin // @[RegSlices.scala 130:31]
      bwd_data_mrkr_req <= io_upStream_bits_mrkr_req;
    end
    if (bwd_ready) begin // @[RegSlices.scala 130:31]
      bwd_data_sdi <= io_upStream_bits_sdi;
    end
    if (bwd_ready) begin // @[RegSlices.scala 130:31]
      bwd_data_qid <= io_upStream_bits_qid;
    end
    if (bwd_ready) begin // @[RegSlices.scala 130:31]
      bwd_data_error <= io_upStream_bits_error;
    end
    if (bwd_ready) begin // @[RegSlices.scala 130:31]
      bwd_data_func <= io_upStream_bits_func;
    end
    if (bwd_ready) begin // @[RegSlices.scala 130:31]
      bwd_data_cidx <= io_upStream_bits_cidx;
    end
    if (bwd_ready) begin // @[RegSlices.scala 130:31]
      bwd_data_port_id <= io_upStream_bits_port_id;
    end
    if (bwd_ready) begin // @[RegSlices.scala 130:31]
      bwd_data_no_dma <= io_upStream_bits_no_dma;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  fwd_valid = _RAND_0[0:0];
  _RAND_1 = {2{`RANDOM}};
  fwd_data_addr = _RAND_1[63:0];
  _RAND_2 = {1{`RANDOM}};
  fwd_data_len = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  fwd_data_eop = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  fwd_data_sop = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  fwd_data_mrkr_req = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  fwd_data_sdi = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  fwd_data_qid = _RAND_7[10:0];
  _RAND_8 = {1{`RANDOM}};
  fwd_data_error = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  fwd_data_func = _RAND_9[7:0];
  _RAND_10 = {1{`RANDOM}};
  fwd_data_cidx = _RAND_10[15:0];
  _RAND_11 = {1{`RANDOM}};
  fwd_data_port_id = _RAND_11[2:0];
  _RAND_12 = {1{`RANDOM}};
  fwd_data_no_dma = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  bwd_ready = _RAND_13[0:0];
  _RAND_14 = {2{`RANDOM}};
  bwd_data_addr = _RAND_14[63:0];
  _RAND_15 = {1{`RANDOM}};
  bwd_data_len = _RAND_15[31:0];
  _RAND_16 = {1{`RANDOM}};
  bwd_data_eop = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  bwd_data_sop = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  bwd_data_mrkr_req = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  bwd_data_sdi = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  bwd_data_qid = _RAND_20[10:0];
  _RAND_21 = {1{`RANDOM}};
  bwd_data_error = _RAND_21[0:0];
  _RAND_22 = {1{`RANDOM}};
  bwd_data_func = _RAND_22[7:0];
  _RAND_23 = {1{`RANDOM}};
  bwd_data_cidx = _RAND_23[15:0];
  _RAND_24 = {1{`RANDOM}};
  bwd_data_port_id = _RAND_24[2:0];
  _RAND_25 = {1{`RANDOM}};
  bwd_data_no_dma = _RAND_25[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module SV_STREAM_FIFO_3(
  input          io_m_clk,
  input          io_s_clk,
  input          io_reset_n,
  input  [127:0] io_in_data,
  input          io_in_valid,
  output         io_in_ready,
  output [127:0] io_out_data,
  output         io_out_valid,
  input          io_out_ready
);
  wire [127:0] meta_m_axis_tdata; // @[Meta.scala 30:26]
  wire [15:0] meta_m_axis_tkeep; // @[Meta.scala 30:26]
  wire  meta_m_axis_tlast; // @[Meta.scala 30:26]
  wire  meta_m_axis_tvalid; // @[Meta.scala 30:26]
  wire [4:0] meta_rd_data_count_axis; // @[Meta.scala 30:26]
  wire  meta_s_axis_tready; // @[Meta.scala 30:26]
  wire [4:0] meta_wr_data_count_axis; // @[Meta.scala 30:26]
  wire  meta_m_aclk; // @[Meta.scala 30:26]
  wire  meta_m_axis_tready; // @[Meta.scala 30:26]
  wire  meta_s_aclk; // @[Meta.scala 30:26]
  wire  meta_s_aresetn; // @[Meta.scala 30:26]
  wire [127:0] meta_s_axis_tdata; // @[Meta.scala 30:26]
  wire  meta_s_axis_tdest; // @[Meta.scala 30:26]
  wire  meta_s_axis_tid; // @[Meta.scala 30:26]
  wire [15:0] meta_s_axis_tkeep; // @[Meta.scala 30:26]
  wire  meta_s_axis_tlast; // @[Meta.scala 30:26]
  wire [15:0] meta_s_axis_tstrb; // @[Meta.scala 30:26]
  wire  meta_s_axis_tuser; // @[Meta.scala 30:26]
  wire  meta_s_axis_tvalid; // @[Meta.scala 30:26]
  xpm_fifo_axis
    #(.RD_DATA_COUNT_WIDTH(5), .CLOCKING_MODE("independent_clock"), .PACKET_FIFO("false"), .USE_ADV_FEATURES("0404"), .TID_WIDTH(1), .TDEST_WIDTH(1), .PROG_EMPTY_THRESH(10), .TUSER_WIDTH(1), .FIFO_DEPTH(16), .SIM_ASSERT_CHK(0), .WR_DATA_COUNT_WIDTH(5), .ECC_MODE("no_ecc"), .FIFO_MEMORY_TYPE("auto"), .PROG_FULL_THRESH(10), .TDATA_WIDTH(128), .RELATED_CLOCKS(0), .CASCADE_HEIGHT(0), .CDC_SYNC_STAGES(2))
    meta ( // @[Meta.scala 30:26]
    .m_axis_tdata(meta_m_axis_tdata),
    .m_axis_tkeep(meta_m_axis_tkeep),
    .m_axis_tlast(meta_m_axis_tlast),
    .m_axis_tvalid(meta_m_axis_tvalid),
    .rd_data_count_axis(meta_rd_data_count_axis),
    .s_axis_tready(meta_s_axis_tready),
    .wr_data_count_axis(meta_wr_data_count_axis),
    .m_aclk(meta_m_aclk),
    .m_axis_tready(meta_m_axis_tready),
    .s_aclk(meta_s_aclk),
    .s_aresetn(meta_s_aresetn),
    .s_axis_tdata(meta_s_axis_tdata),
    .s_axis_tdest(meta_s_axis_tdest),
    .s_axis_tid(meta_s_axis_tid),
    .s_axis_tkeep(meta_s_axis_tkeep),
    .s_axis_tlast(meta_s_axis_tlast),
    .s_axis_tstrb(meta_s_axis_tstrb),
    .s_axis_tuser(meta_s_axis_tuser),
    .s_axis_tvalid(meta_s_axis_tvalid)
  );
  assign io_in_ready = meta_s_axis_tready; // @[Meta.scala 34:41]
  assign io_out_data = meta_m_axis_tdata; // @[Meta.scala 31:41]
  assign io_out_valid = meta_m_axis_tvalid; // @[Meta.scala 32:41]
  assign meta_m_aclk = io_m_clk; // @[Meta.scala 37:49]
  assign meta_m_axis_tready = io_out_ready; // @[Meta.scala 38:41]
  assign meta_s_aclk = io_s_clk; // @[Meta.scala 39:49]
  assign meta_s_aresetn = io_reset_n; // @[Meta.scala 40:49]
  assign meta_s_axis_tdata = io_in_data; // @[Meta.scala 41:41]
  assign meta_s_axis_tdest = 1'h0; // @[Meta.scala 42:41]
  assign meta_s_axis_tid = 1'h0; // @[Meta.scala 43:49]
  assign meta_s_axis_tkeep = 16'hffff; // @[Bitwise.scala 72:12]
  assign meta_s_axis_tlast = 1'h1; // @[Meta.scala 45:41]
  assign meta_s_axis_tstrb = 16'hffff; // @[Bitwise.scala 72:12]
  assign meta_s_axis_tuser = 1'h0; // @[Meta.scala 47:41]
  assign meta_s_axis_tvalid = io_in_valid; // @[Meta.scala 48:41]
endmodule
module XConverter_3(
  input         io_in_clk,
  input         io_out_clk,
  input         io_rstn,
  output        io_in_ready,
  input         io_in_valid,
  input  [63:0] io_in_bits_addr,
  input  [10:0] io_in_bits_qid,
  input         io_in_bits_error,
  input  [7:0]  io_in_bits_func,
  input  [2:0]  io_in_bits_port_id,
  input  [6:0]  io_in_bits_pfch_tag,
  input  [31:0] io_in_bits_len,
  input         io_out_ready,
  output        io_out_valid,
  output [63:0] io_out_bits_addr,
  output [10:0] io_out_bits_qid,
  output        io_out_bits_error,
  output [7:0]  io_out_bits_func,
  output [2:0]  io_out_bits_port_id,
  output [6:0]  io_out_bits_pfch_tag,
  output [31:0] io_out_bits_len,
  output        io_out_ready_0,
  output        io_out_valid_1
);
  wire  fifo_io_m_clk; // @[XConverter.scala 97:34]
  wire  fifo_io_s_clk; // @[XConverter.scala 97:34]
  wire  fifo_io_reset_n; // @[XConverter.scala 97:34]
  wire [127:0] fifo_io_in_data; // @[XConverter.scala 97:34]
  wire  fifo_io_in_valid; // @[XConverter.scala 97:34]
  wire  fifo_io_in_ready; // @[XConverter.scala 97:34]
  wire [127:0] fifo_io_out_data; // @[XConverter.scala 97:34]
  wire  fifo_io_out_valid; // @[XConverter.scala 97:34]
  wire  fifo_io_out_ready; // @[XConverter.scala 97:34]
  wire [125:0] _fifo_io_in_data_T = {io_in_bits_addr,io_in_bits_qid,io_in_bits_error,io_in_bits_func,io_in_bits_port_id,
    io_in_bits_pfch_tag,io_in_bits_len}; // @[XConverter.scala 103:63]
  SV_STREAM_FIFO_3 fifo ( // @[XConverter.scala 97:34]
    .io_m_clk(fifo_io_m_clk),
    .io_s_clk(fifo_io_s_clk),
    .io_reset_n(fifo_io_reset_n),
    .io_in_data(fifo_io_in_data),
    .io_in_valid(fifo_io_in_valid),
    .io_in_ready(fifo_io_in_ready),
    .io_out_data(fifo_io_out_data),
    .io_out_valid(fifo_io_out_valid),
    .io_out_ready(fifo_io_out_ready)
  );
  assign io_in_ready = fifo_io_in_ready; // @[XConverter.scala 105:41]
  assign io_out_valid = fifo_io_out_valid; // @[XConverter.scala 108:41]
  assign io_out_bits_addr = fifo_io_out_data[125:62]; // @[XConverter.scala 107:77]
  assign io_out_bits_qid = fifo_io_out_data[61:51]; // @[XConverter.scala 107:77]
  assign io_out_bits_error = fifo_io_out_data[50]; // @[XConverter.scala 107:77]
  assign io_out_bits_func = fifo_io_out_data[49:42]; // @[XConverter.scala 107:77]
  assign io_out_bits_port_id = fifo_io_out_data[41:39]; // @[XConverter.scala 107:77]
  assign io_out_bits_pfch_tag = fifo_io_out_data[38:32]; // @[XConverter.scala 107:77]
  assign io_out_bits_len = fifo_io_out_data[31:0]; // @[XConverter.scala 107:77]
  assign io_out_ready_0 = io_out_ready;
  assign io_out_valid_1 = io_out_valid;
  assign fifo_io_m_clk = io_out_clk; // @[XConverter.scala 100:41]
  assign fifo_io_s_clk = io_in_clk; // @[XConverter.scala 99:41]
  assign fifo_io_reset_n = io_rstn; // @[XConverter.scala 101:41]
  assign fifo_io_in_data = {{2'd0}, _fifo_io_in_data_T}; // @[XConverter.scala 103:63]
  assign fifo_io_in_valid = io_in_valid; // @[XConverter.scala 104:41]
  assign fifo_io_out_ready = io_out_ready; // @[XConverter.scala 109:41]
endmodule
module RegSlice_3(
  input         clock,
  input         reset,
  output        io_upStream_ready,
  input         io_upStream_valid,
  input  [63:0] io_upStream_bits_addr,
  input  [10:0] io_upStream_bits_qid,
  input         io_upStream_bits_error,
  input  [7:0]  io_upStream_bits_func,
  input  [2:0]  io_upStream_bits_port_id,
  input  [6:0]  io_upStream_bits_pfch_tag,
  input  [31:0] io_upStream_bits_len,
  input         io_downStream_ready,
  output        io_downStream_valid,
  output [63:0] io_downStream_bits_addr,
  output [10:0] io_downStream_bits_qid,
  output        io_downStream_bits_error,
  output [7:0]  io_downStream_bits_func,
  output [2:0]  io_downStream_bits_port_id,
  output [6:0]  io_downStream_bits_pfch_tag,
  output [31:0] io_downStream_bits_len
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [63:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
`endif // RANDOMIZE_REG_INIT
  reg  fwd_valid; // @[RegSlices.scala 112:34]
  reg [63:0] fwd_data_addr; // @[RegSlices.scala 113:30]
  reg [10:0] fwd_data_qid; // @[RegSlices.scala 113:30]
  reg  fwd_data_error; // @[RegSlices.scala 113:30]
  reg [7:0] fwd_data_func; // @[RegSlices.scala 113:30]
  reg [2:0] fwd_data_port_id; // @[RegSlices.scala 113:30]
  reg [6:0] fwd_data_pfch_tag; // @[RegSlices.scala 113:30]
  reg [31:0] fwd_data_len; // @[RegSlices.scala 113:30]
  wire  fwd_ready_s = ~fwd_valid | io_downStream_ready; // @[RegSlices.scala 115:35]
  reg  bwd_ready; // @[RegSlices.scala 123:34]
  reg [63:0] bwd_data_addr; // @[RegSlices.scala 124:30]
  reg [10:0] bwd_data_qid; // @[RegSlices.scala 124:30]
  reg  bwd_data_error; // @[RegSlices.scala 124:30]
  reg [7:0] bwd_data_func; // @[RegSlices.scala 124:30]
  reg [2:0] bwd_data_port_id; // @[RegSlices.scala 124:30]
  reg [6:0] bwd_data_pfch_tag; // @[RegSlices.scala 124:30]
  reg [31:0] bwd_data_len; // @[RegSlices.scala 124:30]
  wire  _fwd_valid_T = io_downStream_ready ? 1'h0 : fwd_valid; // @[RegSlices.scala 121:53]
  wire  bwd_valid_s = ~bwd_ready | io_upStream_valid; // @[RegSlices.scala 126:39]
  wire  _bwd_ready_T = io_upStream_valid ? 1'h0 : bwd_ready; // @[RegSlices.scala 132:53]
  assign io_upStream_ready = bwd_ready; // @[RegSlices.scala 107:31 RegSlices.scala 128:25]
  assign io_downStream_valid = fwd_valid; // @[RegSlices.scala 109:31 RegSlices.scala 116:21]
  assign io_downStream_bits_addr = fwd_data_addr; // @[RegSlices.scala 108:31 RegSlices.scala 117:25]
  assign io_downStream_bits_qid = fwd_data_qid; // @[RegSlices.scala 108:31 RegSlices.scala 117:25]
  assign io_downStream_bits_error = fwd_data_error; // @[RegSlices.scala 108:31 RegSlices.scala 117:25]
  assign io_downStream_bits_func = fwd_data_func; // @[RegSlices.scala 108:31 RegSlices.scala 117:25]
  assign io_downStream_bits_port_id = fwd_data_port_id; // @[RegSlices.scala 108:31 RegSlices.scala 117:25]
  assign io_downStream_bits_pfch_tag = fwd_data_pfch_tag; // @[RegSlices.scala 108:31 RegSlices.scala 117:25]
  assign io_downStream_bits_len = fwd_data_len; // @[RegSlices.scala 108:31 RegSlices.scala 117:25]
  always @(posedge clock) begin
    if (reset) begin // @[RegSlices.scala 112:34]
      fwd_valid <= 1'h0; // @[RegSlices.scala 112:34]
    end else begin
      fwd_valid <= bwd_valid_s | _fwd_valid_T; // @[RegSlices.scala 121:25]
    end
    if (fwd_ready_s) begin // @[RegSlices.scala 119:31]
      if (bwd_ready) begin // @[RegSlices.scala 127:31]
        fwd_data_addr <= io_upStream_bits_addr;
      end else begin
        fwd_data_addr <= bwd_data_addr;
      end
    end
    if (fwd_ready_s) begin // @[RegSlices.scala 119:31]
      if (bwd_ready) begin // @[RegSlices.scala 127:31]
        fwd_data_qid <= io_upStream_bits_qid;
      end else begin
        fwd_data_qid <= bwd_data_qid;
      end
    end
    if (fwd_ready_s) begin // @[RegSlices.scala 119:31]
      if (bwd_ready) begin // @[RegSlices.scala 127:31]
        fwd_data_error <= io_upStream_bits_error;
      end else begin
        fwd_data_error <= bwd_data_error;
      end
    end
    if (fwd_ready_s) begin // @[RegSlices.scala 119:31]
      if (bwd_ready) begin // @[RegSlices.scala 127:31]
        fwd_data_func <= io_upStream_bits_func;
      end else begin
        fwd_data_func <= bwd_data_func;
      end
    end
    if (fwd_ready_s) begin // @[RegSlices.scala 119:31]
      if (bwd_ready) begin // @[RegSlices.scala 127:31]
        fwd_data_port_id <= io_upStream_bits_port_id;
      end else begin
        fwd_data_port_id <= bwd_data_port_id;
      end
    end
    if (fwd_ready_s) begin // @[RegSlices.scala 119:31]
      if (bwd_ready) begin // @[RegSlices.scala 127:31]
        fwd_data_pfch_tag <= io_upStream_bits_pfch_tag;
      end else begin
        fwd_data_pfch_tag <= bwd_data_pfch_tag;
      end
    end
    if (fwd_ready_s) begin // @[RegSlices.scala 119:31]
      if (bwd_ready) begin // @[RegSlices.scala 127:31]
        fwd_data_len <= io_upStream_bits_len;
      end else begin
        fwd_data_len <= bwd_data_len;
      end
    end
    bwd_ready <= reset | (fwd_ready_s | _bwd_ready_T); // @[RegSlices.scala 123:34 RegSlices.scala 123:34 RegSlices.scala 132:25]
    if (bwd_ready) begin // @[RegSlices.scala 130:31]
      bwd_data_addr <= io_upStream_bits_addr;
    end
    if (bwd_ready) begin // @[RegSlices.scala 130:31]
      bwd_data_qid <= io_upStream_bits_qid;
    end
    if (bwd_ready) begin // @[RegSlices.scala 130:31]
      bwd_data_error <= io_upStream_bits_error;
    end
    if (bwd_ready) begin // @[RegSlices.scala 130:31]
      bwd_data_func <= io_upStream_bits_func;
    end
    if (bwd_ready) begin // @[RegSlices.scala 130:31]
      bwd_data_port_id <= io_upStream_bits_port_id;
    end
    if (bwd_ready) begin // @[RegSlices.scala 130:31]
      bwd_data_pfch_tag <= io_upStream_bits_pfch_tag;
    end
    if (bwd_ready) begin // @[RegSlices.scala 130:31]
      bwd_data_len <= io_upStream_bits_len;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  fwd_valid = _RAND_0[0:0];
  _RAND_1 = {2{`RANDOM}};
  fwd_data_addr = _RAND_1[63:0];
  _RAND_2 = {1{`RANDOM}};
  fwd_data_qid = _RAND_2[10:0];
  _RAND_3 = {1{`RANDOM}};
  fwd_data_error = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  fwd_data_func = _RAND_4[7:0];
  _RAND_5 = {1{`RANDOM}};
  fwd_data_port_id = _RAND_5[2:0];
  _RAND_6 = {1{`RANDOM}};
  fwd_data_pfch_tag = _RAND_6[6:0];
  _RAND_7 = {1{`RANDOM}};
  fwd_data_len = _RAND_7[31:0];
  _RAND_8 = {1{`RANDOM}};
  bwd_ready = _RAND_8[0:0];
  _RAND_9 = {2{`RANDOM}};
  bwd_data_addr = _RAND_9[63:0];
  _RAND_10 = {1{`RANDOM}};
  bwd_data_qid = _RAND_10[10:0];
  _RAND_11 = {1{`RANDOM}};
  bwd_data_error = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  bwd_data_func = _RAND_12[7:0];
  _RAND_13 = {1{`RANDOM}};
  bwd_data_port_id = _RAND_13[2:0];
  _RAND_14 = {1{`RANDOM}};
  bwd_data_pfch_tag = _RAND_14[6:0];
  _RAND_15 = {1{`RANDOM}};
  bwd_data_len = _RAND_15[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module CMDBoundaryCheck(
  input         clock,
  input         reset,
  output        io_in_ready,
  input         io_in_valid,
  input  [63:0] io_in_bits_addr,
  input  [10:0] io_in_bits_qid,
  input         io_in_bits_error,
  input  [7:0]  io_in_bits_func,
  input  [2:0]  io_in_bits_port_id,
  input  [6:0]  io_in_bits_pfch_tag,
  input  [31:0] io_in_bits_len,
  input         io_out_ready,
  output        io_out_valid,
  output [63:0] io_out_bits_addr,
  output [10:0] io_out_bits_qid,
  output        io_out_bits_error,
  output [7:0]  io_out_bits_func,
  output [2:0]  io_out_bits_port_id,
  output [6:0]  io_out_bits_pfch_tag,
  output [31:0] io_out_bits_len
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
`endif // RANDOMIZE_REG_INIT
  reg [23:0] offset_addr; // @[CheckSplit.scala 81:34]
  reg [23:0] new_length; // @[CheckSplit.scala 82:33]
  reg [63:0] cmd_addr; // @[CheckSplit.scala 83:31]
  reg [31:0] cmd_len; // @[CheckSplit.scala 84:30]
  reg [63:0] mini_addr; // @[CheckSplit.scala 85:32]
  reg [31:0] mini_len; // @[CheckSplit.scala 86:31]
  reg [10:0] cmd_temp_qid; // @[CheckSplit.scala 87:27]
  reg  cmd_temp_error; // @[CheckSplit.scala 87:27]
  reg [7:0] cmd_temp_func; // @[CheckSplit.scala 87:27]
  reg [2:0] cmd_temp_port_id; // @[CheckSplit.scala 87:27]
  reg [6:0] cmd_temp_pfch_tag; // @[CheckSplit.scala 87:27]
  reg [2:0] state; // @[CheckSplit.scala 90:50]
  wire  _T = 3'h0 == state; // @[Conditional.scala 37:30]
  wire  _T_1 = io_in_ready & io_in_valid; // @[Decoupled.scala 40:37]
  wire [63:0] _offset_addr_T = io_in_bits_addr & 64'h1fffff; // @[CheckSplit.scala 103:92]
  wire [63:0] _new_length_T_2 = 64'h200000 - _offset_addr_T; // @[CheckSplit.scala 105:88]
  wire [63:0] _GEN_9 = _T_1 ? _offset_addr_T : {{40'd0}, offset_addr}; // @[CheckSplit.scala 99:43 CheckSplit.scala 103:73 CheckSplit.scala 81:34]
  wire [63:0] _GEN_11 = _T_1 ? _new_length_T_2 : {{40'd0}, new_length}; // @[CheckSplit.scala 99:43 CheckSplit.scala 105:73 CheckSplit.scala 82:33]
  wire  _T_2 = 3'h1 == state; // @[Conditional.scala 37:30]
  wire [31:0] _GEN_136 = {{8'd0}, offset_addr}; // @[CheckSplit.scala 109:43]
  wire [31:0] _T_4 = _GEN_136 + cmd_len; // @[CheckSplit.scala 109:43]
  wire [63:0] _GEN_137 = {{40'd0}, new_length}; // @[CheckSplit.scala 112:85]
  wire [63:0] _cmd_addr_T_1 = cmd_addr + _GEN_137; // @[CheckSplit.scala 112:85]
  wire [31:0] _GEN_138 = {{8'd0}, new_length}; // @[CheckSplit.scala 113:84]
  wire [31:0] _cmd_len_T_1 = cmd_len - _GEN_138; // @[CheckSplit.scala 113:84]
  wire  _T_6 = 3'h2 == state; // @[Conditional.scala 37:30]
  wire [63:0] _cmd_addr_T_3 = cmd_addr + 64'h200000; // @[CheckSplit.scala 125:85]
  wire [31:0] _cmd_len_T_3 = cmd_len - 32'h200000; // @[CheckSplit.scala 126:84]
  wire [31:0] _GEN_18 = cmd_len > 32'h200000 ? 32'h200000 : cmd_len; // @[CheckSplit.scala 122:52 CheckSplit.scala 124:73 CheckSplit.scala 130:73]
  wire [63:0] _GEN_19 = cmd_len > 32'h200000 ? _cmd_addr_T_3 : cmd_addr; // @[CheckSplit.scala 122:52 CheckSplit.scala 125:73 CheckSplit.scala 83:31]
  wire [31:0] _GEN_20 = cmd_len > 32'h200000 ? _cmd_len_T_3 : cmd_len; // @[CheckSplit.scala 122:52 CheckSplit.scala 126:73 CheckSplit.scala 84:30]
  wire [2:0] _GEN_21 = cmd_len > 32'h200000 ? 3'h3 : 3'h4; // @[CheckSplit.scala 122:52 CheckSplit.scala 127:57 CheckSplit.scala 131:57]
  wire  _T_8 = 3'h3 == state; // @[Conditional.scala 37:30]
  wire  _T_10 = mini_len > 32'h1000; // @[CheckSplit.scala 136:47]
  wire [63:0] _mini_addr_T_1 = mini_addr + 64'h1000; // @[CheckSplit.scala 137:94]
  wire [31:0] _mini_len_T_1 = mini_len - 32'h1000; // @[CheckSplit.scala 138:93]
  wire [63:0] _GEN_22 = mini_len > 32'h1000 ? _mini_addr_T_1 : mini_addr; // @[CheckSplit.scala 136:66 CheckSplit.scala 137:81 CheckSplit.scala 85:32]
  wire [31:0] _GEN_23 = mini_len > 32'h1000 ? _mini_len_T_1 : mini_len; // @[CheckSplit.scala 136:66 CheckSplit.scala 138:81 CheckSplit.scala 86:31]
  wire [31:0] _GEN_25 = mini_len > 32'h1000 ? 32'h1000 : mini_len; // @[CheckSplit.scala 136:66 CheckSplit.scala 141:73 CheckSplit.scala 146:73]
  wire [2:0] _GEN_32 = mini_len > 32'h1000 ? state : 3'h2; // @[CheckSplit.scala 136:66 CheckSplit.scala 90:50 CheckSplit.scala 148:81]
  wire [63:0] _GEN_33 = io_out_ready ? _GEN_22 : mini_addr; // @[CheckSplit.scala 135:51 CheckSplit.scala 85:32]
  wire [31:0] _GEN_34 = io_out_ready ? _GEN_23 : mini_len; // @[CheckSplit.scala 135:51 CheckSplit.scala 86:31]
  wire [31:0] _GEN_36 = io_out_ready ? _GEN_25 : 32'h0; // @[CheckSplit.scala 135:51 CheckSplit.scala 95:65]
  wire [6:0] _GEN_37 = io_out_ready ? cmd_temp_pfch_tag : 7'h0; // @[CheckSplit.scala 135:51 CheckSplit.scala 95:65]
  wire [2:0] _GEN_38 = io_out_ready ? cmd_temp_port_id : 3'h0; // @[CheckSplit.scala 135:51 CheckSplit.scala 95:65]
  wire [7:0] _GEN_39 = io_out_ready ? cmd_temp_func : 8'h0; // @[CheckSplit.scala 135:51 CheckSplit.scala 95:65]
  wire  _GEN_40 = io_out_ready & cmd_temp_error; // @[CheckSplit.scala 135:51 CheckSplit.scala 95:65]
  wire [10:0] _GEN_41 = io_out_ready ? cmd_temp_qid : 11'h0; // @[CheckSplit.scala 135:51 CheckSplit.scala 95:65]
  wire [63:0] _GEN_42 = io_out_ready ? mini_addr : 64'h0; // @[CheckSplit.scala 135:51 CheckSplit.scala 95:65]
  wire [2:0] _GEN_43 = io_out_ready ? _GEN_32 : state; // @[CheckSplit.scala 135:51 CheckSplit.scala 90:50]
  wire  _T_11 = 3'h4 == state; // @[Conditional.scala 37:30]
  wire [2:0] _GEN_54 = _T_10 ? state : 3'h0; // @[CheckSplit.scala 154:66 CheckSplit.scala 90:50 CheckSplit.scala 166:81]
  wire [2:0] _GEN_65 = io_out_ready ? _GEN_54 : state; // @[CheckSplit.scala 153:51 CheckSplit.scala 90:50]
  wire [63:0] _GEN_66 = _T_11 ? _GEN_33 : mini_addr; // @[Conditional.scala 39:67 CheckSplit.scala 85:32]
  wire [31:0] _GEN_67 = _T_11 ? _GEN_34 : mini_len; // @[Conditional.scala 39:67 CheckSplit.scala 86:31]
  wire  _GEN_68 = _T_11 & io_out_ready; // @[Conditional.scala 39:67 CheckSplit.scala 94:57]
  wire [31:0] _GEN_69 = _T_11 ? _GEN_36 : 32'h0; // @[Conditional.scala 39:67 CheckSplit.scala 95:65]
  wire [6:0] _GEN_70 = _T_11 ? _GEN_37 : 7'h0; // @[Conditional.scala 39:67 CheckSplit.scala 95:65]
  wire [2:0] _GEN_71 = _T_11 ? _GEN_38 : 3'h0; // @[Conditional.scala 39:67 CheckSplit.scala 95:65]
  wire [7:0] _GEN_72 = _T_11 ? _GEN_39 : 8'h0; // @[Conditional.scala 39:67 CheckSplit.scala 95:65]
  wire  _GEN_73 = _T_11 & _GEN_40; // @[Conditional.scala 39:67 CheckSplit.scala 95:65]
  wire [10:0] _GEN_74 = _T_11 ? _GEN_41 : 11'h0; // @[Conditional.scala 39:67 CheckSplit.scala 95:65]
  wire [63:0] _GEN_75 = _T_11 ? _GEN_42 : 64'h0; // @[Conditional.scala 39:67 CheckSplit.scala 95:65]
  wire [2:0] _GEN_76 = _T_11 ? _GEN_65 : state; // @[Conditional.scala 39:67 CheckSplit.scala 90:50]
  wire [63:0] _GEN_77 = _T_8 ? _GEN_33 : _GEN_66; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_78 = _T_8 ? _GEN_34 : _GEN_67; // @[Conditional.scala 39:67]
  wire  _GEN_79 = _T_8 ? io_out_ready : _GEN_68; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_80 = _T_8 ? _GEN_36 : _GEN_69; // @[Conditional.scala 39:67]
  wire [6:0] _GEN_81 = _T_8 ? _GEN_37 : _GEN_70; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_82 = _T_8 ? _GEN_38 : _GEN_71; // @[Conditional.scala 39:67]
  wire [7:0] _GEN_83 = _T_8 ? _GEN_39 : _GEN_72; // @[Conditional.scala 39:67]
  wire  _GEN_84 = _T_8 ? _GEN_40 : _GEN_73; // @[Conditional.scala 39:67]
  wire [10:0] _GEN_85 = _T_8 ? _GEN_41 : _GEN_74; // @[Conditional.scala 39:67]
  wire [63:0] _GEN_86 = _T_8 ? _GEN_42 : _GEN_75; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_87 = _T_8 ? _GEN_43 : _GEN_76; // @[Conditional.scala 39:67]
  wire  _GEN_93 = _T_6 ? 1'h0 : _GEN_79; // @[Conditional.scala 39:67 CheckSplit.scala 94:57]
  wire [31:0] _GEN_94 = _T_6 ? 32'h0 : _GEN_80; // @[Conditional.scala 39:67 CheckSplit.scala 95:65]
  wire [6:0] _GEN_95 = _T_6 ? 7'h0 : _GEN_81; // @[Conditional.scala 39:67 CheckSplit.scala 95:65]
  wire [2:0] _GEN_96 = _T_6 ? 3'h0 : _GEN_82; // @[Conditional.scala 39:67 CheckSplit.scala 95:65]
  wire [7:0] _GEN_97 = _T_6 ? 8'h0 : _GEN_83; // @[Conditional.scala 39:67 CheckSplit.scala 95:65]
  wire  _GEN_98 = _T_6 ? 1'h0 : _GEN_84; // @[Conditional.scala 39:67 CheckSplit.scala 95:65]
  wire [10:0] _GEN_99 = _T_6 ? 11'h0 : _GEN_85; // @[Conditional.scala 39:67 CheckSplit.scala 95:65]
  wire [63:0] _GEN_100 = _T_6 ? 64'h0 : _GEN_86; // @[Conditional.scala 39:67 CheckSplit.scala 95:65]
  wire  _GEN_106 = _T_2 ? 1'h0 : _GEN_93; // @[Conditional.scala 39:67 CheckSplit.scala 94:57]
  wire [31:0] _GEN_107 = _T_2 ? 32'h0 : _GEN_94; // @[Conditional.scala 39:67 CheckSplit.scala 95:65]
  wire [6:0] _GEN_108 = _T_2 ? 7'h0 : _GEN_95; // @[Conditional.scala 39:67 CheckSplit.scala 95:65]
  wire [2:0] _GEN_109 = _T_2 ? 3'h0 : _GEN_96; // @[Conditional.scala 39:67 CheckSplit.scala 95:65]
  wire [7:0] _GEN_110 = _T_2 ? 8'h0 : _GEN_97; // @[Conditional.scala 39:67 CheckSplit.scala 95:65]
  wire  _GEN_111 = _T_2 ? 1'h0 : _GEN_98; // @[Conditional.scala 39:67 CheckSplit.scala 95:65]
  wire [10:0] _GEN_112 = _T_2 ? 11'h0 : _GEN_99; // @[Conditional.scala 39:67 CheckSplit.scala 95:65]
  wire [63:0] _GEN_113 = _T_2 ? 64'h0 : _GEN_100; // @[Conditional.scala 39:67 CheckSplit.scala 95:65]
  wire [63:0] _GEN_123 = _T ? _GEN_9 : {{40'd0}, offset_addr}; // @[Conditional.scala 40:58 CheckSplit.scala 81:34]
  wire [63:0] _GEN_125 = _T ? _GEN_11 : {{40'd0}, new_length}; // @[Conditional.scala 40:58 CheckSplit.scala 82:33]
  assign io_in_ready = state == 3'h0; // @[CheckSplit.scala 92:75]
  assign io_out_valid = _T ? 1'h0 : _GEN_106; // @[Conditional.scala 40:58 CheckSplit.scala 94:57]
  assign io_out_bits_addr = _T ? 64'h0 : _GEN_113; // @[Conditional.scala 40:58 CheckSplit.scala 95:65]
  assign io_out_bits_qid = _T ? 11'h0 : _GEN_112; // @[Conditional.scala 40:58 CheckSplit.scala 95:65]
  assign io_out_bits_error = _T ? 1'h0 : _GEN_111; // @[Conditional.scala 40:58 CheckSplit.scala 95:65]
  assign io_out_bits_func = _T ? 8'h0 : _GEN_110; // @[Conditional.scala 40:58 CheckSplit.scala 95:65]
  assign io_out_bits_port_id = _T ? 3'h0 : _GEN_109; // @[Conditional.scala 40:58 CheckSplit.scala 95:65]
  assign io_out_bits_pfch_tag = _T ? 7'h0 : _GEN_108; // @[Conditional.scala 40:58 CheckSplit.scala 95:65]
  assign io_out_bits_len = _T ? 32'h0 : _GEN_107; // @[Conditional.scala 40:58 CheckSplit.scala 95:65]
  always @(posedge clock) begin
    if (reset) begin // @[CheckSplit.scala 81:34]
      offset_addr <= 24'h0; // @[CheckSplit.scala 81:34]
    end else begin
      offset_addr <= _GEN_123[23:0];
    end
    if (reset) begin // @[CheckSplit.scala 82:33]
      new_length <= 24'h0; // @[CheckSplit.scala 82:33]
    end else begin
      new_length <= _GEN_125[23:0];
    end
    if (reset) begin // @[CheckSplit.scala 83:31]
      cmd_addr <= 64'h0; // @[CheckSplit.scala 83:31]
    end else if (_T) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[CheckSplit.scala 99:43]
        cmd_addr <= io_in_bits_addr; // @[CheckSplit.scala 100:73]
      end
    end else if (_T_2) begin // @[Conditional.scala 39:67]
      if (_T_4 > 32'h200000) begin // @[CheckSplit.scala 109:68]
        cmd_addr <= _cmd_addr_T_1; // @[CheckSplit.scala 112:73]
      end
    end else if (_T_6) begin // @[Conditional.scala 39:67]
      cmd_addr <= _GEN_19;
    end
    if (reset) begin // @[CheckSplit.scala 84:30]
      cmd_len <= 32'h0; // @[CheckSplit.scala 84:30]
    end else if (_T) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[CheckSplit.scala 99:43]
        cmd_len <= io_in_bits_len; // @[CheckSplit.scala 101:73]
      end
    end else if (_T_2) begin // @[Conditional.scala 39:67]
      if (_T_4 > 32'h200000) begin // @[CheckSplit.scala 109:68]
        cmd_len <= _cmd_len_T_1; // @[CheckSplit.scala 113:73]
      end
    end else if (_T_6) begin // @[Conditional.scala 39:67]
      cmd_len <= _GEN_20;
    end
    if (reset) begin // @[CheckSplit.scala 85:32]
      mini_addr <= 64'h0; // @[CheckSplit.scala 85:32]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_2) begin // @[Conditional.scala 39:67]
        mini_addr <= cmd_addr;
      end else if (_T_6) begin // @[Conditional.scala 39:67]
        mini_addr <= cmd_addr;
      end else begin
        mini_addr <= _GEN_77;
      end
    end
    if (reset) begin // @[CheckSplit.scala 86:31]
      mini_len <= 32'h0; // @[CheckSplit.scala 86:31]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_2) begin // @[Conditional.scala 39:67]
        if (_T_4 > 32'h200000) begin // @[CheckSplit.scala 109:68]
          mini_len <= {{8'd0}, new_length}; // @[CheckSplit.scala 111:73]
        end else begin
          mini_len <= cmd_len; // @[CheckSplit.scala 117:73]
        end
      end else if (_T_6) begin // @[Conditional.scala 39:67]
        mini_len <= _GEN_18;
      end else begin
        mini_len <= _GEN_78;
      end
    end
    if (_T) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[CheckSplit.scala 99:43]
        cmd_temp_qid <= io_in_bits_qid; // @[CheckSplit.scala 102:73]
      end
    end
    if (_T) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[CheckSplit.scala 99:43]
        cmd_temp_error <= io_in_bits_error; // @[CheckSplit.scala 102:73]
      end
    end
    if (_T) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[CheckSplit.scala 99:43]
        cmd_temp_func <= io_in_bits_func; // @[CheckSplit.scala 102:73]
      end
    end
    if (_T) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[CheckSplit.scala 99:43]
        cmd_temp_port_id <= io_in_bits_port_id; // @[CheckSplit.scala 102:73]
      end
    end
    if (_T) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[CheckSplit.scala 99:43]
        cmd_temp_pfch_tag <= io_in_bits_pfch_tag; // @[CheckSplit.scala 102:73]
      end
    end
    if (reset) begin // @[CheckSplit.scala 90:50]
      state <= 3'h0; // @[CheckSplit.scala 90:50]
    end else if (_T) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[CheckSplit.scala 99:43]
        state <= 3'h1; // @[CheckSplit.scala 104:41]
      end
    end else if (_T_2) begin // @[Conditional.scala 39:67]
      if (_T_4 > 32'h200000) begin // @[CheckSplit.scala 109:68]
        state <= 3'h3; // @[CheckSplit.scala 114:57]
      end else begin
        state <= 3'h4; // @[CheckSplit.scala 118:57]
      end
    end else if (_T_6) begin // @[Conditional.scala 39:67]
      state <= _GEN_21;
    end else begin
      state <= _GEN_87;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  offset_addr = _RAND_0[23:0];
  _RAND_1 = {1{`RANDOM}};
  new_length = _RAND_1[23:0];
  _RAND_2 = {2{`RANDOM}};
  cmd_addr = _RAND_2[63:0];
  _RAND_3 = {1{`RANDOM}};
  cmd_len = _RAND_3[31:0];
  _RAND_4 = {2{`RANDOM}};
  mini_addr = _RAND_4[63:0];
  _RAND_5 = {1{`RANDOM}};
  mini_len = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  cmd_temp_qid = _RAND_6[10:0];
  _RAND_7 = {1{`RANDOM}};
  cmd_temp_error = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  cmd_temp_func = _RAND_8[7:0];
  _RAND_9 = {1{`RANDOM}};
  cmd_temp_port_id = _RAND_9[2:0];
  _RAND_10 = {1{`RANDOM}};
  cmd_temp_pfch_tag = _RAND_10[6:0];
  _RAND_11 = {1{`RANDOM}};
  state = _RAND_11[2:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module CMDBoundaryCheck_1(
  input         clock,
  input         reset,
  output        io_in_ready,
  input         io_in_valid,
  input  [63:0] io_in_bits_addr,
  input  [31:0] io_in_bits_len,
  input         io_in_bits_eop,
  input         io_in_bits_sop,
  input         io_in_bits_mrkr_req,
  input         io_in_bits_sdi,
  input  [10:0] io_in_bits_qid,
  input         io_in_bits_error,
  input  [7:0]  io_in_bits_func,
  input  [15:0] io_in_bits_cidx,
  input  [2:0]  io_in_bits_port_id,
  input         io_in_bits_no_dma,
  input         io_out_ready,
  output        io_out_valid,
  output [63:0] io_out_bits_addr,
  output [31:0] io_out_bits_len,
  output        io_out_bits_eop,
  output        io_out_bits_sop,
  output        io_out_bits_mrkr_req,
  output        io_out_bits_sdi,
  output [10:0] io_out_bits_qid,
  output        io_out_bits_error,
  output [7:0]  io_out_bits_func,
  output [15:0] io_out_bits_cidx,
  output [2:0]  io_out_bits_port_id,
  output        io_out_bits_no_dma
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
`endif // RANDOMIZE_REG_INIT
  reg [23:0] offset_addr; // @[CheckSplit.scala 81:34]
  reg [23:0] new_length; // @[CheckSplit.scala 82:33]
  reg [63:0] cmd_addr; // @[CheckSplit.scala 83:31]
  reg [31:0] cmd_len; // @[CheckSplit.scala 84:30]
  reg [63:0] mini_addr; // @[CheckSplit.scala 85:32]
  reg [31:0] mini_len; // @[CheckSplit.scala 86:31]
  reg  cmd_temp_eop; // @[CheckSplit.scala 87:27]
  reg  cmd_temp_sop; // @[CheckSplit.scala 87:27]
  reg  cmd_temp_mrkr_req; // @[CheckSplit.scala 87:27]
  reg  cmd_temp_sdi; // @[CheckSplit.scala 87:27]
  reg [10:0] cmd_temp_qid; // @[CheckSplit.scala 87:27]
  reg  cmd_temp_error; // @[CheckSplit.scala 87:27]
  reg [7:0] cmd_temp_func; // @[CheckSplit.scala 87:27]
  reg [15:0] cmd_temp_cidx; // @[CheckSplit.scala 87:27]
  reg [2:0] cmd_temp_port_id; // @[CheckSplit.scala 87:27]
  reg  cmd_temp_no_dma; // @[CheckSplit.scala 87:27]
  reg [2:0] state; // @[CheckSplit.scala 90:50]
  wire  _T = 3'h0 == state; // @[Conditional.scala 37:30]
  wire  _T_1 = io_in_ready & io_in_valid; // @[Decoupled.scala 40:37]
  wire [63:0] _offset_addr_T = io_in_bits_addr & 64'h1fffff; // @[CheckSplit.scala 103:92]
  wire [63:0] _new_length_T_2 = 64'h200000 - _offset_addr_T; // @[CheckSplit.scala 105:88]
  wire [63:0] _GEN_14 = _T_1 ? _offset_addr_T : {{40'd0}, offset_addr}; // @[CheckSplit.scala 99:43 CheckSplit.scala 103:73 CheckSplit.scala 81:34]
  wire [63:0] _GEN_16 = _T_1 ? _new_length_T_2 : {{40'd0}, new_length}; // @[CheckSplit.scala 99:43 CheckSplit.scala 105:73 CheckSplit.scala 82:33]
  wire  _T_2 = 3'h1 == state; // @[Conditional.scala 37:30]
  wire [31:0] _GEN_191 = {{8'd0}, offset_addr}; // @[CheckSplit.scala 109:43]
  wire [31:0] _T_4 = _GEN_191 + cmd_len; // @[CheckSplit.scala 109:43]
  wire [63:0] _GEN_192 = {{40'd0}, new_length}; // @[CheckSplit.scala 112:85]
  wire [63:0] _cmd_addr_T_1 = cmd_addr + _GEN_192; // @[CheckSplit.scala 112:85]
  wire [31:0] _GEN_193 = {{8'd0}, new_length}; // @[CheckSplit.scala 113:84]
  wire [31:0] _cmd_len_T_1 = cmd_len - _GEN_193; // @[CheckSplit.scala 113:84]
  wire  _T_6 = 3'h2 == state; // @[Conditional.scala 37:30]
  wire [63:0] _cmd_addr_T_3 = cmd_addr + 64'h200000; // @[CheckSplit.scala 125:85]
  wire [31:0] _cmd_len_T_3 = cmd_len - 32'h200000; // @[CheckSplit.scala 126:84]
  wire [31:0] _GEN_23 = cmd_len > 32'h200000 ? 32'h200000 : cmd_len; // @[CheckSplit.scala 122:52 CheckSplit.scala 124:73 CheckSplit.scala 130:73]
  wire [63:0] _GEN_24 = cmd_len > 32'h200000 ? _cmd_addr_T_3 : cmd_addr; // @[CheckSplit.scala 122:52 CheckSplit.scala 125:73 CheckSplit.scala 83:31]
  wire [31:0] _GEN_25 = cmd_len > 32'h200000 ? _cmd_len_T_3 : cmd_len; // @[CheckSplit.scala 122:52 CheckSplit.scala 126:73 CheckSplit.scala 84:30]
  wire [2:0] _GEN_26 = cmd_len > 32'h200000 ? 3'h3 : 3'h4; // @[CheckSplit.scala 122:52 CheckSplit.scala 127:57 CheckSplit.scala 131:57]
  wire  _T_8 = 3'h3 == state; // @[Conditional.scala 37:30]
  wire  _T_10 = mini_len > 32'h8000; // @[CheckSplit.scala 136:47]
  wire [63:0] _mini_addr_T_1 = mini_addr + 64'h8000; // @[CheckSplit.scala 137:94]
  wire [31:0] _mini_len_T_1 = mini_len - 32'h8000; // @[CheckSplit.scala 138:93]
  wire [63:0] _GEN_27 = mini_len > 32'h8000 ? _mini_addr_T_1 : mini_addr; // @[CheckSplit.scala 136:66 CheckSplit.scala 137:81 CheckSplit.scala 85:32]
  wire [31:0] _GEN_28 = mini_len > 32'h8000 ? _mini_len_T_1 : mini_len; // @[CheckSplit.scala 136:66 CheckSplit.scala 138:81 CheckSplit.scala 86:31]
  wire [31:0] _GEN_40 = mini_len > 32'h8000 ? 32'h8000 : mini_len; // @[CheckSplit.scala 136:66 CheckSplit.scala 141:73 CheckSplit.scala 146:73]
  wire [2:0] _GEN_42 = mini_len > 32'h8000 ? state : 3'h2; // @[CheckSplit.scala 136:66 CheckSplit.scala 90:50 CheckSplit.scala 148:81]
  wire [63:0] _GEN_43 = io_out_ready ? _GEN_27 : mini_addr; // @[CheckSplit.scala 135:51 CheckSplit.scala 85:32]
  wire [31:0] _GEN_44 = io_out_ready ? _GEN_28 : mini_len; // @[CheckSplit.scala 135:51 CheckSplit.scala 86:31]
  wire  _GEN_46 = io_out_ready & cmd_temp_no_dma; // @[CheckSplit.scala 135:51 CheckSplit.scala 95:65]
  wire [2:0] _GEN_47 = io_out_ready ? cmd_temp_port_id : 3'h0; // @[CheckSplit.scala 135:51 CheckSplit.scala 95:65]
  wire [15:0] _GEN_48 = io_out_ready ? cmd_temp_cidx : 16'h0; // @[CheckSplit.scala 135:51 CheckSplit.scala 95:65]
  wire [7:0] _GEN_49 = io_out_ready ? cmd_temp_func : 8'h0; // @[CheckSplit.scala 135:51 CheckSplit.scala 95:65]
  wire  _GEN_50 = io_out_ready & cmd_temp_error; // @[CheckSplit.scala 135:51 CheckSplit.scala 95:65]
  wire [10:0] _GEN_51 = io_out_ready ? cmd_temp_qid : 11'h0; // @[CheckSplit.scala 135:51 CheckSplit.scala 95:65]
  wire  _GEN_52 = io_out_ready & cmd_temp_sdi; // @[CheckSplit.scala 135:51 CheckSplit.scala 95:65]
  wire  _GEN_53 = io_out_ready & cmd_temp_mrkr_req; // @[CheckSplit.scala 135:51 CheckSplit.scala 95:65]
  wire  _GEN_54 = io_out_ready & cmd_temp_sop; // @[CheckSplit.scala 135:51 CheckSplit.scala 95:65]
  wire  _GEN_55 = io_out_ready & cmd_temp_eop; // @[CheckSplit.scala 135:51 CheckSplit.scala 95:65]
  wire [31:0] _GEN_56 = io_out_ready ? _GEN_40 : 32'h0; // @[CheckSplit.scala 135:51 CheckSplit.scala 95:65]
  wire [63:0] _GEN_57 = io_out_ready ? mini_addr : 64'h0; // @[CheckSplit.scala 135:51 CheckSplit.scala 95:65]
  wire [2:0] _GEN_58 = io_out_ready ? _GEN_42 : state; // @[CheckSplit.scala 135:51 CheckSplit.scala 90:50]
  wire  _T_11 = 3'h4 == state; // @[Conditional.scala 37:30]
  wire [2:0] _GEN_74 = _T_10 ? state : 3'h0; // @[CheckSplit.scala 154:66 CheckSplit.scala 90:50 CheckSplit.scala 166:81]
  wire [2:0] _GEN_90 = io_out_ready ? _GEN_74 : state; // @[CheckSplit.scala 153:51 CheckSplit.scala 90:50]
  wire [63:0] _GEN_91 = _T_11 ? _GEN_43 : mini_addr; // @[Conditional.scala 39:67 CheckSplit.scala 85:32]
  wire [31:0] _GEN_92 = _T_11 ? _GEN_44 : mini_len; // @[Conditional.scala 39:67 CheckSplit.scala 86:31]
  wire  _GEN_93 = _T_11 & io_out_ready; // @[Conditional.scala 39:67 CheckSplit.scala 94:57]
  wire  _GEN_94 = _T_11 & _GEN_46; // @[Conditional.scala 39:67 CheckSplit.scala 95:65]
  wire [2:0] _GEN_95 = _T_11 ? _GEN_47 : 3'h0; // @[Conditional.scala 39:67 CheckSplit.scala 95:65]
  wire [15:0] _GEN_96 = _T_11 ? _GEN_48 : 16'h0; // @[Conditional.scala 39:67 CheckSplit.scala 95:65]
  wire [7:0] _GEN_97 = _T_11 ? _GEN_49 : 8'h0; // @[Conditional.scala 39:67 CheckSplit.scala 95:65]
  wire  _GEN_98 = _T_11 & _GEN_50; // @[Conditional.scala 39:67 CheckSplit.scala 95:65]
  wire [10:0] _GEN_99 = _T_11 ? _GEN_51 : 11'h0; // @[Conditional.scala 39:67 CheckSplit.scala 95:65]
  wire  _GEN_100 = _T_11 & _GEN_52; // @[Conditional.scala 39:67 CheckSplit.scala 95:65]
  wire  _GEN_101 = _T_11 & _GEN_53; // @[Conditional.scala 39:67 CheckSplit.scala 95:65]
  wire  _GEN_102 = _T_11 & _GEN_54; // @[Conditional.scala 39:67 CheckSplit.scala 95:65]
  wire  _GEN_103 = _T_11 & _GEN_55; // @[Conditional.scala 39:67 CheckSplit.scala 95:65]
  wire [31:0] _GEN_104 = _T_11 ? _GEN_56 : 32'h0; // @[Conditional.scala 39:67 CheckSplit.scala 95:65]
  wire [63:0] _GEN_105 = _T_11 ? _GEN_57 : 64'h0; // @[Conditional.scala 39:67 CheckSplit.scala 95:65]
  wire [2:0] _GEN_106 = _T_11 ? _GEN_90 : state; // @[Conditional.scala 39:67 CheckSplit.scala 90:50]
  wire [63:0] _GEN_107 = _T_8 ? _GEN_43 : _GEN_91; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_108 = _T_8 ? _GEN_44 : _GEN_92; // @[Conditional.scala 39:67]
  wire  _GEN_109 = _T_8 ? io_out_ready : _GEN_93; // @[Conditional.scala 39:67]
  wire  _GEN_110 = _T_8 ? _GEN_46 : _GEN_94; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_111 = _T_8 ? _GEN_47 : _GEN_95; // @[Conditional.scala 39:67]
  wire [15:0] _GEN_112 = _T_8 ? _GEN_48 : _GEN_96; // @[Conditional.scala 39:67]
  wire [7:0] _GEN_113 = _T_8 ? _GEN_49 : _GEN_97; // @[Conditional.scala 39:67]
  wire  _GEN_114 = _T_8 ? _GEN_50 : _GEN_98; // @[Conditional.scala 39:67]
  wire [10:0] _GEN_115 = _T_8 ? _GEN_51 : _GEN_99; // @[Conditional.scala 39:67]
  wire  _GEN_116 = _T_8 ? _GEN_52 : _GEN_100; // @[Conditional.scala 39:67]
  wire  _GEN_117 = _T_8 ? _GEN_53 : _GEN_101; // @[Conditional.scala 39:67]
  wire  _GEN_118 = _T_8 ? _GEN_54 : _GEN_102; // @[Conditional.scala 39:67]
  wire  _GEN_119 = _T_8 ? _GEN_55 : _GEN_103; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_120 = _T_8 ? _GEN_56 : _GEN_104; // @[Conditional.scala 39:67]
  wire [63:0] _GEN_121 = _T_8 ? _GEN_57 : _GEN_105; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_122 = _T_8 ? _GEN_58 : _GEN_106; // @[Conditional.scala 39:67]
  wire  _GEN_128 = _T_6 ? 1'h0 : _GEN_109; // @[Conditional.scala 39:67 CheckSplit.scala 94:57]
  wire  _GEN_129 = _T_6 ? 1'h0 : _GEN_110; // @[Conditional.scala 39:67 CheckSplit.scala 95:65]
  wire [2:0] _GEN_130 = _T_6 ? 3'h0 : _GEN_111; // @[Conditional.scala 39:67 CheckSplit.scala 95:65]
  wire [15:0] _GEN_131 = _T_6 ? 16'h0 : _GEN_112; // @[Conditional.scala 39:67 CheckSplit.scala 95:65]
  wire [7:0] _GEN_132 = _T_6 ? 8'h0 : _GEN_113; // @[Conditional.scala 39:67 CheckSplit.scala 95:65]
  wire  _GEN_133 = _T_6 ? 1'h0 : _GEN_114; // @[Conditional.scala 39:67 CheckSplit.scala 95:65]
  wire [10:0] _GEN_134 = _T_6 ? 11'h0 : _GEN_115; // @[Conditional.scala 39:67 CheckSplit.scala 95:65]
  wire  _GEN_135 = _T_6 ? 1'h0 : _GEN_116; // @[Conditional.scala 39:67 CheckSplit.scala 95:65]
  wire  _GEN_136 = _T_6 ? 1'h0 : _GEN_117; // @[Conditional.scala 39:67 CheckSplit.scala 95:65]
  wire  _GEN_137 = _T_6 ? 1'h0 : _GEN_118; // @[Conditional.scala 39:67 CheckSplit.scala 95:65]
  wire  _GEN_138 = _T_6 ? 1'h0 : _GEN_119; // @[Conditional.scala 39:67 CheckSplit.scala 95:65]
  wire [31:0] _GEN_139 = _T_6 ? 32'h0 : _GEN_120; // @[Conditional.scala 39:67 CheckSplit.scala 95:65]
  wire [63:0] _GEN_140 = _T_6 ? 64'h0 : _GEN_121; // @[Conditional.scala 39:67 CheckSplit.scala 95:65]
  wire  _GEN_146 = _T_2 ? 1'h0 : _GEN_128; // @[Conditional.scala 39:67 CheckSplit.scala 94:57]
  wire  _GEN_147 = _T_2 ? 1'h0 : _GEN_129; // @[Conditional.scala 39:67 CheckSplit.scala 95:65]
  wire [2:0] _GEN_148 = _T_2 ? 3'h0 : _GEN_130; // @[Conditional.scala 39:67 CheckSplit.scala 95:65]
  wire [15:0] _GEN_149 = _T_2 ? 16'h0 : _GEN_131; // @[Conditional.scala 39:67 CheckSplit.scala 95:65]
  wire [7:0] _GEN_150 = _T_2 ? 8'h0 : _GEN_132; // @[Conditional.scala 39:67 CheckSplit.scala 95:65]
  wire  _GEN_151 = _T_2 ? 1'h0 : _GEN_133; // @[Conditional.scala 39:67 CheckSplit.scala 95:65]
  wire [10:0] _GEN_152 = _T_2 ? 11'h0 : _GEN_134; // @[Conditional.scala 39:67 CheckSplit.scala 95:65]
  wire  _GEN_153 = _T_2 ? 1'h0 : _GEN_135; // @[Conditional.scala 39:67 CheckSplit.scala 95:65]
  wire  _GEN_154 = _T_2 ? 1'h0 : _GEN_136; // @[Conditional.scala 39:67 CheckSplit.scala 95:65]
  wire  _GEN_155 = _T_2 ? 1'h0 : _GEN_137; // @[Conditional.scala 39:67 CheckSplit.scala 95:65]
  wire  _GEN_156 = _T_2 ? 1'h0 : _GEN_138; // @[Conditional.scala 39:67 CheckSplit.scala 95:65]
  wire [31:0] _GEN_157 = _T_2 ? 32'h0 : _GEN_139; // @[Conditional.scala 39:67 CheckSplit.scala 95:65]
  wire [63:0] _GEN_158 = _T_2 ? 64'h0 : _GEN_140; // @[Conditional.scala 39:67 CheckSplit.scala 95:65]
  wire [63:0] _GEN_173 = _T ? _GEN_14 : {{40'd0}, offset_addr}; // @[Conditional.scala 40:58 CheckSplit.scala 81:34]
  wire [63:0] _GEN_175 = _T ? _GEN_16 : {{40'd0}, new_length}; // @[Conditional.scala 40:58 CheckSplit.scala 82:33]
  assign io_in_ready = state == 3'h0; // @[CheckSplit.scala 92:75]
  assign io_out_valid = _T ? 1'h0 : _GEN_146; // @[Conditional.scala 40:58 CheckSplit.scala 94:57]
  assign io_out_bits_addr = _T ? 64'h0 : _GEN_158; // @[Conditional.scala 40:58 CheckSplit.scala 95:65]
  assign io_out_bits_len = _T ? 32'h0 : _GEN_157; // @[Conditional.scala 40:58 CheckSplit.scala 95:65]
  assign io_out_bits_eop = _T ? 1'h0 : _GEN_156; // @[Conditional.scala 40:58 CheckSplit.scala 95:65]
  assign io_out_bits_sop = _T ? 1'h0 : _GEN_155; // @[Conditional.scala 40:58 CheckSplit.scala 95:65]
  assign io_out_bits_mrkr_req = _T ? 1'h0 : _GEN_154; // @[Conditional.scala 40:58 CheckSplit.scala 95:65]
  assign io_out_bits_sdi = _T ? 1'h0 : _GEN_153; // @[Conditional.scala 40:58 CheckSplit.scala 95:65]
  assign io_out_bits_qid = _T ? 11'h0 : _GEN_152; // @[Conditional.scala 40:58 CheckSplit.scala 95:65]
  assign io_out_bits_error = _T ? 1'h0 : _GEN_151; // @[Conditional.scala 40:58 CheckSplit.scala 95:65]
  assign io_out_bits_func = _T ? 8'h0 : _GEN_150; // @[Conditional.scala 40:58 CheckSplit.scala 95:65]
  assign io_out_bits_cidx = _T ? 16'h0 : _GEN_149; // @[Conditional.scala 40:58 CheckSplit.scala 95:65]
  assign io_out_bits_port_id = _T ? 3'h0 : _GEN_148; // @[Conditional.scala 40:58 CheckSplit.scala 95:65]
  assign io_out_bits_no_dma = _T ? 1'h0 : _GEN_147; // @[Conditional.scala 40:58 CheckSplit.scala 95:65]
  always @(posedge clock) begin
    if (reset) begin // @[CheckSplit.scala 81:34]
      offset_addr <= 24'h0; // @[CheckSplit.scala 81:34]
    end else begin
      offset_addr <= _GEN_173[23:0];
    end
    if (reset) begin // @[CheckSplit.scala 82:33]
      new_length <= 24'h0; // @[CheckSplit.scala 82:33]
    end else begin
      new_length <= _GEN_175[23:0];
    end
    if (reset) begin // @[CheckSplit.scala 83:31]
      cmd_addr <= 64'h0; // @[CheckSplit.scala 83:31]
    end else if (_T) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[CheckSplit.scala 99:43]
        cmd_addr <= io_in_bits_addr; // @[CheckSplit.scala 100:73]
      end
    end else if (_T_2) begin // @[Conditional.scala 39:67]
      if (_T_4 > 32'h200000) begin // @[CheckSplit.scala 109:68]
        cmd_addr <= _cmd_addr_T_1; // @[CheckSplit.scala 112:73]
      end
    end else if (_T_6) begin // @[Conditional.scala 39:67]
      cmd_addr <= _GEN_24;
    end
    if (reset) begin // @[CheckSplit.scala 84:30]
      cmd_len <= 32'h0; // @[CheckSplit.scala 84:30]
    end else if (_T) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[CheckSplit.scala 99:43]
        cmd_len <= io_in_bits_len; // @[CheckSplit.scala 101:73]
      end
    end else if (_T_2) begin // @[Conditional.scala 39:67]
      if (_T_4 > 32'h200000) begin // @[CheckSplit.scala 109:68]
        cmd_len <= _cmd_len_T_1; // @[CheckSplit.scala 113:73]
      end
    end else if (_T_6) begin // @[Conditional.scala 39:67]
      cmd_len <= _GEN_25;
    end
    if (reset) begin // @[CheckSplit.scala 85:32]
      mini_addr <= 64'h0; // @[CheckSplit.scala 85:32]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_2) begin // @[Conditional.scala 39:67]
        mini_addr <= cmd_addr;
      end else if (_T_6) begin // @[Conditional.scala 39:67]
        mini_addr <= cmd_addr;
      end else begin
        mini_addr <= _GEN_107;
      end
    end
    if (reset) begin // @[CheckSplit.scala 86:31]
      mini_len <= 32'h0; // @[CheckSplit.scala 86:31]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_2) begin // @[Conditional.scala 39:67]
        if (_T_4 > 32'h200000) begin // @[CheckSplit.scala 109:68]
          mini_len <= {{8'd0}, new_length}; // @[CheckSplit.scala 111:73]
        end else begin
          mini_len <= cmd_len; // @[CheckSplit.scala 117:73]
        end
      end else if (_T_6) begin // @[Conditional.scala 39:67]
        mini_len <= _GEN_23;
      end else begin
        mini_len <= _GEN_108;
      end
    end
    if (_T) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[CheckSplit.scala 99:43]
        cmd_temp_eop <= io_in_bits_eop; // @[CheckSplit.scala 102:73]
      end
    end
    if (_T) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[CheckSplit.scala 99:43]
        cmd_temp_sop <= io_in_bits_sop; // @[CheckSplit.scala 102:73]
      end
    end
    if (_T) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[CheckSplit.scala 99:43]
        cmd_temp_mrkr_req <= io_in_bits_mrkr_req; // @[CheckSplit.scala 102:73]
      end
    end
    if (_T) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[CheckSplit.scala 99:43]
        cmd_temp_sdi <= io_in_bits_sdi; // @[CheckSplit.scala 102:73]
      end
    end
    if (_T) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[CheckSplit.scala 99:43]
        cmd_temp_qid <= io_in_bits_qid; // @[CheckSplit.scala 102:73]
      end
    end
    if (_T) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[CheckSplit.scala 99:43]
        cmd_temp_error <= io_in_bits_error; // @[CheckSplit.scala 102:73]
      end
    end
    if (_T) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[CheckSplit.scala 99:43]
        cmd_temp_func <= io_in_bits_func; // @[CheckSplit.scala 102:73]
      end
    end
    if (_T) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[CheckSplit.scala 99:43]
        cmd_temp_cidx <= io_in_bits_cidx; // @[CheckSplit.scala 102:73]
      end
    end
    if (_T) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[CheckSplit.scala 99:43]
        cmd_temp_port_id <= io_in_bits_port_id; // @[CheckSplit.scala 102:73]
      end
    end
    if (_T) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[CheckSplit.scala 99:43]
        cmd_temp_no_dma <= io_in_bits_no_dma; // @[CheckSplit.scala 102:73]
      end
    end
    if (reset) begin // @[CheckSplit.scala 90:50]
      state <= 3'h0; // @[CheckSplit.scala 90:50]
    end else if (_T) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[CheckSplit.scala 99:43]
        state <= 3'h1; // @[CheckSplit.scala 104:41]
      end
    end else if (_T_2) begin // @[Conditional.scala 39:67]
      if (_T_4 > 32'h200000) begin // @[CheckSplit.scala 109:68]
        state <= 3'h3; // @[CheckSplit.scala 114:57]
      end else begin
        state <= 3'h4; // @[CheckSplit.scala 118:57]
      end
    end else if (_T_6) begin // @[Conditional.scala 39:67]
      state <= _GEN_26;
    end else begin
      state <= _GEN_122;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  offset_addr = _RAND_0[23:0];
  _RAND_1 = {1{`RANDOM}};
  new_length = _RAND_1[23:0];
  _RAND_2 = {2{`RANDOM}};
  cmd_addr = _RAND_2[63:0];
  _RAND_3 = {1{`RANDOM}};
  cmd_len = _RAND_3[31:0];
  _RAND_4 = {2{`RANDOM}};
  mini_addr = _RAND_4[63:0];
  _RAND_5 = {1{`RANDOM}};
  mini_len = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  cmd_temp_eop = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  cmd_temp_sop = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  cmd_temp_mrkr_req = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  cmd_temp_sdi = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  cmd_temp_qid = _RAND_10[10:0];
  _RAND_11 = {1{`RANDOM}};
  cmd_temp_error = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  cmd_temp_func = _RAND_12[7:0];
  _RAND_13 = {1{`RANDOM}};
  cmd_temp_cidx = _RAND_13[15:0];
  _RAND_14 = {1{`RANDOM}};
  cmd_temp_port_id = _RAND_14[2:0];
  _RAND_15 = {1{`RANDOM}};
  cmd_temp_no_dma = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  state = _RAND_16[2:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module XRam(
  input         clock,
  input         reset,
  input  [12:0] io_addr_a,
  input  [12:0] io_addr_b,
  input         io_wr_en_a,
  input  [63:0] io_data_in_a,
  output [63:0] io_data_out_a,
  output [63:0] io_data_out_b
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [63:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [63:0] _RAND_16;
  reg [63:0] _RAND_17;
`endif // RANDOMIZE_REG_INIT
  wire [63:0] ram_douta; // @[XRam.scala 136:33]
  wire [63:0] ram_doutb; // @[XRam.scala 136:33]
  wire [12:0] ram_addra; // @[XRam.scala 136:33]
  wire [12:0] ram_addrb; // @[XRam.scala 136:33]
  wire  ram_clka; // @[XRam.scala 136:33]
  wire  ram_clkb; // @[XRam.scala 136:33]
  wire [63:0] ram_dina; // @[XRam.scala 136:33]
  wire [63:0] ram_dinb; // @[XRam.scala 136:33]
  wire  ram_ena; // @[XRam.scala 136:33]
  wire  ram_enb; // @[XRam.scala 136:33]
  wire  ram_injectdbiterra; // @[XRam.scala 136:33]
  wire  ram_injectdbiterrb; // @[XRam.scala 136:33]
  wire  ram_injectsbiterra; // @[XRam.scala 136:33]
  wire  ram_injectsbiterrb; // @[XRam.scala 136:33]
  wire  ram_regcea; // @[XRam.scala 136:33]
  wire  ram_regceb; // @[XRam.scala 136:33]
  wire  ram_rsta; // @[XRam.scala 136:33]
  wire  ram_rstb; // @[XRam.scala 136:33]
  wire  ram_sleep; // @[XRam.scala 136:33]
  wire [7:0] ram_wea; // @[XRam.scala 136:33]
  wire [7:0] ram_web; // @[XRam.scala 136:33]
  wire [7:0] wr_en_a = io_wr_en_a ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  reg  usr_rst_delay_r; // @[Reg.scala 15:16]
  reg  usr_rst_delay_r_1; // @[Reg.scala 15:16]
  reg  usr_rst_delay_r_2; // @[Reg.scala 15:16]
  reg  usr_rst_delay; // @[Reg.scala 15:16]
  reg [12:0] reset_addr; // @[XRam.scala 141:54]
  wire [12:0] _reset_addr_T_1 = reset_addr + 13'h1; // @[XRam.scala 144:70]
  reg [12:0] r; // @[Reg.scala 15:16]
  reg [12:0] r_1; // @[Reg.scala 15:16]
  reg [12:0] REG; // @[XRam.scala 165:74]
  reg  REG_1; // @[XRam.scala 165:95]
  reg [63:0] io_data_out_b_REG; // @[XRam.scala 166:75]
  reg [12:0] r_2; // @[Reg.scala 15:16]
  reg [12:0] r_3; // @[Reg.scala 15:16]
  reg [12:0] r_4; // @[Reg.scala 15:16]
  reg [12:0] r_5; // @[Reg.scala 15:16]
  reg  r_6; // @[Reg.scala 15:16]
  reg  r_7; // @[Reg.scala 15:16]
  reg [63:0] io_data_out_b_r; // @[Reg.scala 15:16]
  reg [63:0] io_data_out_b_r_1; // @[Reg.scala 15:16]
  wire [63:0] _io_data_out_b_WIRE = ram_doutb; // @[XRam.scala 170:89 XRam.scala 170:89]
  wire [63:0] _GEN_15 = r_3 == r_5 & r_7 ? io_data_out_b_r_1 : _io_data_out_b_WIRE; // @[XRam.scala 167:130 XRam.scala 168:65 XRam.scala 170:65]
  xpm_memory_tdpram
    #(.USE_EMBEDDED_CONSTRAINT(0), .CLOCKING_MODE("common_clock"), .WRITE_DATA_WIDTH_B(64), .READ_LATENCY_B(2), .ADDR_WIDTH_A(13), .READ_DATA_WIDTH_A(64), .RST_MODE_B("SYNC"), .WAKEUP_TIME("disable_sleep"), .MEMORY_INIT_FILE("none"), .READ_LATENCY_A(2), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_A(64), .AUTO_SLEEP_TIME(0), .WRITE_MODE_A("no_change"), .MEMORY_PRIMITIVE("auto"), .USE_MEM_INIT(1), .MEMORY_INIT_PARAM(""), .SIM_ASSERT_CHK(0), .ECC_MODE("no_ecc"), .READ_RESET_VALUE_A("0"), .BYTE_WRITE_WIDTH_A(8), .MEMORY_OPTIMIZATION("true"), .MESSAGE_CONTROL(0), .WRITE_MODE_B("no_change"), .READ_DATA_WIDTH_B(64), .ADDR_WIDTH_B(13), .CASCADE_HEIGHT(0), .READ_RESET_VALUE_B("0"), .BYTE_WRITE_WIDTH_B(8), .MEMORY_SIZE(524288))
    ram ( // @[XRam.scala 136:33]
    .douta(ram_douta),
    .doutb(ram_doutb),
    .addra(ram_addra),
    .addrb(ram_addrb),
    .clka(ram_clka),
    .clkb(ram_clkb),
    .dina(ram_dina),
    .dinb(ram_dinb),
    .ena(ram_ena),
    .enb(ram_enb),
    .injectdbiterra(ram_injectdbiterra),
    .injectdbiterrb(ram_injectdbiterrb),
    .injectsbiterra(ram_injectsbiterra),
    .injectsbiterrb(ram_injectsbiterrb),
    .regcea(ram_regcea),
    .regceb(ram_regceb),
    .rsta(ram_rsta),
    .rstb(ram_rstb),
    .sleep(ram_sleep),
    .wea(ram_wea),
    .web(ram_web)
  );
  assign io_data_out_a = ram_douta; // @[XRam.scala 175:73 XRam.scala 175:73]
  assign io_data_out_b = r_1 == REG & REG_1 ? io_data_out_b_REG : _GEN_15; // @[XRam.scala 165:108 XRam.scala 166:65]
  assign ram_addra = usr_rst_delay ? reset_addr : io_addr_a; // @[XRam.scala 178:55]
  assign ram_addrb = io_addr_b; // @[XRam.scala 179:49]
  assign ram_clka = clock; // @[XRam.scala 181:57]
  assign ram_clkb = clock; // @[XRam.scala 182:57]
  assign ram_dina = usr_rst_delay ? 64'h0 : io_data_in_a; // @[XRam.scala 184:63]
  assign ram_dinb = 64'h0; // @[XRam.scala 185:57]
  assign ram_ena = 1'h1; // @[XRam.scala 187:57]
  assign ram_enb = 1'h1; // @[XRam.scala 188:57]
  assign ram_injectdbiterra = 1'h0; // @[XRam.scala 190:41]
  assign ram_injectdbiterrb = 1'h0; // @[XRam.scala 191:41]
  assign ram_injectsbiterra = 1'h0; // @[XRam.scala 193:41]
  assign ram_injectsbiterrb = 1'h0; // @[XRam.scala 194:41]
  assign ram_regcea = 1'h1; // @[XRam.scala 196:49]
  assign ram_regceb = 1'h1; // @[XRam.scala 197:49]
  assign ram_rsta = 1'h0; // @[XRam.scala 199:57]
  assign ram_rstb = 1'h0; // @[XRam.scala 200:57]
  assign ram_sleep = 1'h0; // @[XRam.scala 202:49]
  assign ram_wea = usr_rst_delay ? 8'hff : wr_en_a; // @[XRam.scala 206:63]
  assign ram_web = 8'h0; // @[XRam.scala 208:57]
  always @(posedge clock) begin
    usr_rst_delay_r <= reset; // @[Reg.scala 16:19 Reg.scala 16:23 Reg.scala 15:16]
    usr_rst_delay_r_1 <= usr_rst_delay_r; // @[Reg.scala 16:19 Reg.scala 16:23 Reg.scala 15:16]
    usr_rst_delay_r_2 <= usr_rst_delay_r_1; // @[Reg.scala 16:19 Reg.scala 16:23 Reg.scala 15:16]
    usr_rst_delay <= usr_rst_delay_r_2; // @[Reg.scala 16:19 Reg.scala 16:23 Reg.scala 15:16]
    if (usr_rst_delay) begin // @[XRam.scala 143:45]
      reset_addr <= _reset_addr_T_1; // @[XRam.scala 144:57]
    end else begin
      reset_addr <= 13'h0; // @[XRam.scala 146:57]
    end
    r <= io_addr_b; // @[Reg.scala 16:19 Reg.scala 16:23 Reg.scala 15:16]
    r_1 <= r; // @[Reg.scala 16:19 Reg.scala 16:23 Reg.scala 15:16]
    REG <= io_addr_a; // @[XRam.scala 165:74]
    REG_1 <= io_wr_en_a; // @[XRam.scala 165:95]
    io_data_out_b_REG <= io_data_in_a; // @[XRam.scala 166:75]
    r_2 <= io_addr_b; // @[Reg.scala 16:19 Reg.scala 16:23 Reg.scala 15:16]
    r_3 <= r_2; // @[Reg.scala 16:19 Reg.scala 16:23 Reg.scala 15:16]
    r_4 <= io_addr_a; // @[Reg.scala 16:19 Reg.scala 16:23 Reg.scala 15:16]
    r_5 <= r_4; // @[Reg.scala 16:19 Reg.scala 16:23 Reg.scala 15:16]
    r_6 <= io_wr_en_a; // @[Reg.scala 16:19 Reg.scala 16:23 Reg.scala 15:16]
    r_7 <= r_6; // @[Reg.scala 16:19 Reg.scala 16:23 Reg.scala 15:16]
    io_data_out_b_r <= io_data_in_a; // @[Reg.scala 16:19 Reg.scala 16:23 Reg.scala 15:16]
    io_data_out_b_r_1 <= io_data_out_b_r; // @[Reg.scala 16:19 Reg.scala 16:23 Reg.scala 15:16]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  usr_rst_delay_r = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  usr_rst_delay_r_1 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  usr_rst_delay_r_2 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  usr_rst_delay = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  reset_addr = _RAND_4[12:0];
  _RAND_5 = {1{`RANDOM}};
  r = _RAND_5[12:0];
  _RAND_6 = {1{`RANDOM}};
  r_1 = _RAND_6[12:0];
  _RAND_7 = {1{`RANDOM}};
  REG = _RAND_7[12:0];
  _RAND_8 = {1{`RANDOM}};
  REG_1 = _RAND_8[0:0];
  _RAND_9 = {2{`RANDOM}};
  io_data_out_b_REG = _RAND_9[63:0];
  _RAND_10 = {1{`RANDOM}};
  r_2 = _RAND_10[12:0];
  _RAND_11 = {1{`RANDOM}};
  r_3 = _RAND_11[12:0];
  _RAND_12 = {1{`RANDOM}};
  r_4 = _RAND_12[12:0];
  _RAND_13 = {1{`RANDOM}};
  r_5 = _RAND_13[12:0];
  _RAND_14 = {1{`RANDOM}};
  r_6 = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  r_7 = _RAND_15[0:0];
  _RAND_16 = {2{`RANDOM}};
  io_data_out_b_r = _RAND_16[63:0];
  _RAND_17 = {2{`RANDOM}};
  io_data_out_b_r_1 = _RAND_17[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Queue(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input  [63:0] io_enq_bits_addr,
  input  [31:0] io_enq_bits_len,
  input         io_enq_bits_eop,
  input         io_enq_bits_sop,
  input         io_enq_bits_mrkr_req,
  input         io_enq_bits_sdi,
  input  [10:0] io_enq_bits_qid,
  input         io_enq_bits_error,
  input  [7:0]  io_enq_bits_func,
  input  [15:0] io_enq_bits_cidx,
  input  [2:0]  io_enq_bits_port_id,
  input         io_enq_bits_no_dma,
  input         io_deq_ready,
  output        io_deq_valid,
  output [63:0] io_deq_bits_addr,
  output [31:0] io_deq_bits_len,
  output        io_deq_bits_eop,
  output        io_deq_bits_sop,
  output        io_deq_bits_mrkr_req,
  output        io_deq_bits_sdi,
  output [10:0] io_deq_bits_qid,
  output        io_deq_bits_error,
  output [7:0]  io_deq_bits_func,
  output [15:0] io_deq_bits_cidx,
  output [2:0]  io_deq_bits_port_id,
  output        io_deq_bits_no_dma,
  output [3:0]  io_count
);
`ifdef RANDOMIZE_GARBAGE_ASSIGN
  reg [63:0] _RAND_1;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_23;
`endif // RANDOMIZE_GARBAGE_ASSIGN
`ifdef RANDOMIZE_MEM_INIT
  reg [63:0] _RAND_0;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_22;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
`endif // RANDOMIZE_REG_INIT
  reg [63:0] ram_addr [0:9]; // @[Decoupled.scala 218:16]
  wire [63:0] ram_addr_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16]
  wire [3:0] ram_addr_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16]
  wire [63:0] ram_addr_MPORT_data; // @[Decoupled.scala 218:16]
  wire [3:0] ram_addr_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_addr_MPORT_mask; // @[Decoupled.scala 218:16]
  wire  ram_addr_MPORT_en; // @[Decoupled.scala 218:16]
  reg [31:0] ram_len [0:9]; // @[Decoupled.scala 218:16]
  wire [31:0] ram_len_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16]
  wire [3:0] ram_len_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16]
  wire [31:0] ram_len_MPORT_data; // @[Decoupled.scala 218:16]
  wire [3:0] ram_len_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_len_MPORT_mask; // @[Decoupled.scala 218:16]
  wire  ram_len_MPORT_en; // @[Decoupled.scala 218:16]
  reg  ram_eop [0:9]; // @[Decoupled.scala 218:16]
  wire  ram_eop_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16]
  wire [3:0] ram_eop_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_eop_MPORT_data; // @[Decoupled.scala 218:16]
  wire [3:0] ram_eop_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_eop_MPORT_mask; // @[Decoupled.scala 218:16]
  wire  ram_eop_MPORT_en; // @[Decoupled.scala 218:16]
  reg  ram_sop [0:9]; // @[Decoupled.scala 218:16]
  wire  ram_sop_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16]
  wire [3:0] ram_sop_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_sop_MPORT_data; // @[Decoupled.scala 218:16]
  wire [3:0] ram_sop_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_sop_MPORT_mask; // @[Decoupled.scala 218:16]
  wire  ram_sop_MPORT_en; // @[Decoupled.scala 218:16]
  reg  ram_mrkr_req [0:9]; // @[Decoupled.scala 218:16]
  wire  ram_mrkr_req_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16]
  wire [3:0] ram_mrkr_req_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_mrkr_req_MPORT_data; // @[Decoupled.scala 218:16]
  wire [3:0] ram_mrkr_req_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_mrkr_req_MPORT_mask; // @[Decoupled.scala 218:16]
  wire  ram_mrkr_req_MPORT_en; // @[Decoupled.scala 218:16]
  reg  ram_sdi [0:9]; // @[Decoupled.scala 218:16]
  wire  ram_sdi_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16]
  wire [3:0] ram_sdi_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_sdi_MPORT_data; // @[Decoupled.scala 218:16]
  wire [3:0] ram_sdi_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_sdi_MPORT_mask; // @[Decoupled.scala 218:16]
  wire  ram_sdi_MPORT_en; // @[Decoupled.scala 218:16]
  reg [10:0] ram_qid [0:9]; // @[Decoupled.scala 218:16]
  wire [10:0] ram_qid_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16]
  wire [3:0] ram_qid_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16]
  wire [10:0] ram_qid_MPORT_data; // @[Decoupled.scala 218:16]
  wire [3:0] ram_qid_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_qid_MPORT_mask; // @[Decoupled.scala 218:16]
  wire  ram_qid_MPORT_en; // @[Decoupled.scala 218:16]
  reg  ram_error [0:9]; // @[Decoupled.scala 218:16]
  wire  ram_error_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16]
  wire [3:0] ram_error_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_error_MPORT_data; // @[Decoupled.scala 218:16]
  wire [3:0] ram_error_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_error_MPORT_mask; // @[Decoupled.scala 218:16]
  wire  ram_error_MPORT_en; // @[Decoupled.scala 218:16]
  reg [7:0] ram_func [0:9]; // @[Decoupled.scala 218:16]
  wire [7:0] ram_func_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16]
  wire [3:0] ram_func_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16]
  wire [7:0] ram_func_MPORT_data; // @[Decoupled.scala 218:16]
  wire [3:0] ram_func_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_func_MPORT_mask; // @[Decoupled.scala 218:16]
  wire  ram_func_MPORT_en; // @[Decoupled.scala 218:16]
  reg [15:0] ram_cidx [0:9]; // @[Decoupled.scala 218:16]
  wire [15:0] ram_cidx_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16]
  wire [3:0] ram_cidx_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16]
  wire [15:0] ram_cidx_MPORT_data; // @[Decoupled.scala 218:16]
  wire [3:0] ram_cidx_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_cidx_MPORT_mask; // @[Decoupled.scala 218:16]
  wire  ram_cidx_MPORT_en; // @[Decoupled.scala 218:16]
  reg [2:0] ram_port_id [0:9]; // @[Decoupled.scala 218:16]
  wire [2:0] ram_port_id_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16]
  wire [3:0] ram_port_id_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16]
  wire [2:0] ram_port_id_MPORT_data; // @[Decoupled.scala 218:16]
  wire [3:0] ram_port_id_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_port_id_MPORT_mask; // @[Decoupled.scala 218:16]
  wire  ram_port_id_MPORT_en; // @[Decoupled.scala 218:16]
  reg  ram_no_dma [0:9]; // @[Decoupled.scala 218:16]
  wire  ram_no_dma_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16]
  wire [3:0] ram_no_dma_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_no_dma_MPORT_data; // @[Decoupled.scala 218:16]
  wire [3:0] ram_no_dma_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_no_dma_MPORT_mask; // @[Decoupled.scala 218:16]
  wire  ram_no_dma_MPORT_en; // @[Decoupled.scala 218:16]
  reg [3:0] enq_ptr_value; // @[Counter.scala 60:40]
  reg [3:0] deq_ptr_value; // @[Counter.scala 60:40]
  reg  maybe_full; // @[Decoupled.scala 221:27]
  wire  ptr_match = enq_ptr_value == deq_ptr_value; // @[Decoupled.scala 223:33]
  wire  empty = ptr_match & ~maybe_full; // @[Decoupled.scala 224:25]
  wire  full = ptr_match & maybe_full; // @[Decoupled.scala 225:24]
  wire  do_enq = io_enq_ready & io_enq_valid; // @[Decoupled.scala 40:37]
  wire  do_deq = io_deq_ready & io_deq_valid; // @[Decoupled.scala 40:37]
  wire  wrap = enq_ptr_value == 4'h9; // @[Counter.scala 72:24]
  wire [3:0] _value_T_1 = enq_ptr_value + 4'h1; // @[Counter.scala 76:24]
  wire  wrap_1 = deq_ptr_value == 4'h9; // @[Counter.scala 72:24]
  wire [3:0] _value_T_3 = deq_ptr_value + 4'h1; // @[Counter.scala 76:24]
  wire [3:0] ptr_diff = enq_ptr_value - deq_ptr_value; // @[Decoupled.scala 257:32]
  wire [3:0] _io_count_T = maybe_full ? 4'ha : 4'h0; // @[Decoupled.scala 262:24]
  wire [3:0] _io_count_T_3 = 4'ha + ptr_diff; // @[Decoupled.scala 265:38]
  wire [3:0] _io_count_T_4 = deq_ptr_value > enq_ptr_value ? _io_count_T_3 : ptr_diff; // @[Decoupled.scala 264:24]
  assign ram_addr_io_deq_bits_MPORT_addr = deq_ptr_value;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign ram_addr_io_deq_bits_MPORT_data = ram_addr[ram_addr_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  `else
  assign ram_addr_io_deq_bits_MPORT_data = ram_addr_io_deq_bits_MPORT_addr >= 4'ha ? _RAND_1[63:0] :
    ram_addr[ram_addr_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign ram_addr_MPORT_data = io_enq_bits_addr;
  assign ram_addr_MPORT_addr = enq_ptr_value;
  assign ram_addr_MPORT_mask = 1'h1;
  assign ram_addr_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_len_io_deq_bits_MPORT_addr = deq_ptr_value;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign ram_len_io_deq_bits_MPORT_data = ram_len[ram_len_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  `else
  assign ram_len_io_deq_bits_MPORT_data = ram_len_io_deq_bits_MPORT_addr >= 4'ha ? _RAND_3[31:0] :
    ram_len[ram_len_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign ram_len_MPORT_data = io_enq_bits_len;
  assign ram_len_MPORT_addr = enq_ptr_value;
  assign ram_len_MPORT_mask = 1'h1;
  assign ram_len_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_eop_io_deq_bits_MPORT_addr = deq_ptr_value;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign ram_eop_io_deq_bits_MPORT_data = ram_eop[ram_eop_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  `else
  assign ram_eop_io_deq_bits_MPORT_data = ram_eop_io_deq_bits_MPORT_addr >= 4'ha ? _RAND_5[0:0] :
    ram_eop[ram_eop_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign ram_eop_MPORT_data = io_enq_bits_eop;
  assign ram_eop_MPORT_addr = enq_ptr_value;
  assign ram_eop_MPORT_mask = 1'h1;
  assign ram_eop_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_sop_io_deq_bits_MPORT_addr = deq_ptr_value;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign ram_sop_io_deq_bits_MPORT_data = ram_sop[ram_sop_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  `else
  assign ram_sop_io_deq_bits_MPORT_data = ram_sop_io_deq_bits_MPORT_addr >= 4'ha ? _RAND_7[0:0] :
    ram_sop[ram_sop_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign ram_sop_MPORT_data = io_enq_bits_sop;
  assign ram_sop_MPORT_addr = enq_ptr_value;
  assign ram_sop_MPORT_mask = 1'h1;
  assign ram_sop_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_mrkr_req_io_deq_bits_MPORT_addr = deq_ptr_value;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign ram_mrkr_req_io_deq_bits_MPORT_data = ram_mrkr_req[ram_mrkr_req_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  `else
  assign ram_mrkr_req_io_deq_bits_MPORT_data = ram_mrkr_req_io_deq_bits_MPORT_addr >= 4'ha ? _RAND_9[0:0] :
    ram_mrkr_req[ram_mrkr_req_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign ram_mrkr_req_MPORT_data = io_enq_bits_mrkr_req;
  assign ram_mrkr_req_MPORT_addr = enq_ptr_value;
  assign ram_mrkr_req_MPORT_mask = 1'h1;
  assign ram_mrkr_req_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_sdi_io_deq_bits_MPORT_addr = deq_ptr_value;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign ram_sdi_io_deq_bits_MPORT_data = ram_sdi[ram_sdi_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  `else
  assign ram_sdi_io_deq_bits_MPORT_data = ram_sdi_io_deq_bits_MPORT_addr >= 4'ha ? _RAND_11[0:0] :
    ram_sdi[ram_sdi_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign ram_sdi_MPORT_data = io_enq_bits_sdi;
  assign ram_sdi_MPORT_addr = enq_ptr_value;
  assign ram_sdi_MPORT_mask = 1'h1;
  assign ram_sdi_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_qid_io_deq_bits_MPORT_addr = deq_ptr_value;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign ram_qid_io_deq_bits_MPORT_data = ram_qid[ram_qid_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  `else
  assign ram_qid_io_deq_bits_MPORT_data = ram_qid_io_deq_bits_MPORT_addr >= 4'ha ? _RAND_13[10:0] :
    ram_qid[ram_qid_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign ram_qid_MPORT_data = io_enq_bits_qid;
  assign ram_qid_MPORT_addr = enq_ptr_value;
  assign ram_qid_MPORT_mask = 1'h1;
  assign ram_qid_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_error_io_deq_bits_MPORT_addr = deq_ptr_value;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign ram_error_io_deq_bits_MPORT_data = ram_error[ram_error_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  `else
  assign ram_error_io_deq_bits_MPORT_data = ram_error_io_deq_bits_MPORT_addr >= 4'ha ? _RAND_15[0:0] :
    ram_error[ram_error_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign ram_error_MPORT_data = io_enq_bits_error;
  assign ram_error_MPORT_addr = enq_ptr_value;
  assign ram_error_MPORT_mask = 1'h1;
  assign ram_error_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_func_io_deq_bits_MPORT_addr = deq_ptr_value;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign ram_func_io_deq_bits_MPORT_data = ram_func[ram_func_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  `else
  assign ram_func_io_deq_bits_MPORT_data = ram_func_io_deq_bits_MPORT_addr >= 4'ha ? _RAND_17[7:0] :
    ram_func[ram_func_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign ram_func_MPORT_data = io_enq_bits_func;
  assign ram_func_MPORT_addr = enq_ptr_value;
  assign ram_func_MPORT_mask = 1'h1;
  assign ram_func_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_cidx_io_deq_bits_MPORT_addr = deq_ptr_value;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign ram_cidx_io_deq_bits_MPORT_data = ram_cidx[ram_cidx_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  `else
  assign ram_cidx_io_deq_bits_MPORT_data = ram_cidx_io_deq_bits_MPORT_addr >= 4'ha ? _RAND_19[15:0] :
    ram_cidx[ram_cidx_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign ram_cidx_MPORT_data = io_enq_bits_cidx;
  assign ram_cidx_MPORT_addr = enq_ptr_value;
  assign ram_cidx_MPORT_mask = 1'h1;
  assign ram_cidx_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_port_id_io_deq_bits_MPORT_addr = deq_ptr_value;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign ram_port_id_io_deq_bits_MPORT_data = ram_port_id[ram_port_id_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  `else
  assign ram_port_id_io_deq_bits_MPORT_data = ram_port_id_io_deq_bits_MPORT_addr >= 4'ha ? _RAND_21[2:0] :
    ram_port_id[ram_port_id_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign ram_port_id_MPORT_data = io_enq_bits_port_id;
  assign ram_port_id_MPORT_addr = enq_ptr_value;
  assign ram_port_id_MPORT_mask = 1'h1;
  assign ram_port_id_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_no_dma_io_deq_bits_MPORT_addr = deq_ptr_value;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign ram_no_dma_io_deq_bits_MPORT_data = ram_no_dma[ram_no_dma_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  `else
  assign ram_no_dma_io_deq_bits_MPORT_data = ram_no_dma_io_deq_bits_MPORT_addr >= 4'ha ? _RAND_23[0:0] :
    ram_no_dma[ram_no_dma_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign ram_no_dma_MPORT_data = io_enq_bits_no_dma;
  assign ram_no_dma_MPORT_addr = enq_ptr_value;
  assign ram_no_dma_MPORT_mask = 1'h1;
  assign ram_no_dma_MPORT_en = io_enq_ready & io_enq_valid;
  assign io_enq_ready = ~full; // @[Decoupled.scala 241:19]
  assign io_deq_valid = ~empty; // @[Decoupled.scala 240:19]
  assign io_deq_bits_addr = ram_addr_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15]
  assign io_deq_bits_len = ram_len_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15]
  assign io_deq_bits_eop = ram_eop_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15]
  assign io_deq_bits_sop = ram_sop_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15]
  assign io_deq_bits_mrkr_req = ram_mrkr_req_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15]
  assign io_deq_bits_sdi = ram_sdi_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15]
  assign io_deq_bits_qid = ram_qid_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15]
  assign io_deq_bits_error = ram_error_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15]
  assign io_deq_bits_func = ram_func_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15]
  assign io_deq_bits_cidx = ram_cidx_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15]
  assign io_deq_bits_port_id = ram_port_id_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15]
  assign io_deq_bits_no_dma = ram_no_dma_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15]
  assign io_count = ptr_match ? _io_count_T : _io_count_T_4; // @[Decoupled.scala 261:20]
  always @(posedge clock) begin
    if(ram_addr_MPORT_en & ram_addr_MPORT_mask) begin
      ram_addr[ram_addr_MPORT_addr] <= ram_addr_MPORT_data; // @[Decoupled.scala 218:16]
    end
    if(ram_len_MPORT_en & ram_len_MPORT_mask) begin
      ram_len[ram_len_MPORT_addr] <= ram_len_MPORT_data; // @[Decoupled.scala 218:16]
    end
    if(ram_eop_MPORT_en & ram_eop_MPORT_mask) begin
      ram_eop[ram_eop_MPORT_addr] <= ram_eop_MPORT_data; // @[Decoupled.scala 218:16]
    end
    if(ram_sop_MPORT_en & ram_sop_MPORT_mask) begin
      ram_sop[ram_sop_MPORT_addr] <= ram_sop_MPORT_data; // @[Decoupled.scala 218:16]
    end
    if(ram_mrkr_req_MPORT_en & ram_mrkr_req_MPORT_mask) begin
      ram_mrkr_req[ram_mrkr_req_MPORT_addr] <= ram_mrkr_req_MPORT_data; // @[Decoupled.scala 218:16]
    end
    if(ram_sdi_MPORT_en & ram_sdi_MPORT_mask) begin
      ram_sdi[ram_sdi_MPORT_addr] <= ram_sdi_MPORT_data; // @[Decoupled.scala 218:16]
    end
    if(ram_qid_MPORT_en & ram_qid_MPORT_mask) begin
      ram_qid[ram_qid_MPORT_addr] <= ram_qid_MPORT_data; // @[Decoupled.scala 218:16]
    end
    if(ram_error_MPORT_en & ram_error_MPORT_mask) begin
      ram_error[ram_error_MPORT_addr] <= ram_error_MPORT_data; // @[Decoupled.scala 218:16]
    end
    if(ram_func_MPORT_en & ram_func_MPORT_mask) begin
      ram_func[ram_func_MPORT_addr] <= ram_func_MPORT_data; // @[Decoupled.scala 218:16]
    end
    if(ram_cidx_MPORT_en & ram_cidx_MPORT_mask) begin
      ram_cidx[ram_cidx_MPORT_addr] <= ram_cidx_MPORT_data; // @[Decoupled.scala 218:16]
    end
    if(ram_port_id_MPORT_en & ram_port_id_MPORT_mask) begin
      ram_port_id[ram_port_id_MPORT_addr] <= ram_port_id_MPORT_data; // @[Decoupled.scala 218:16]
    end
    if(ram_no_dma_MPORT_en & ram_no_dma_MPORT_mask) begin
      ram_no_dma[ram_no_dma_MPORT_addr] <= ram_no_dma_MPORT_data; // @[Decoupled.scala 218:16]
    end
    if (reset) begin // @[Counter.scala 60:40]
      enq_ptr_value <= 4'h0; // @[Counter.scala 60:40]
    end else if (do_enq) begin // @[Decoupled.scala 229:17]
      if (wrap) begin // @[Counter.scala 86:20]
        enq_ptr_value <= 4'h0; // @[Counter.scala 86:28]
      end else begin
        enq_ptr_value <= _value_T_1; // @[Counter.scala 76:15]
      end
    end
    if (reset) begin // @[Counter.scala 60:40]
      deq_ptr_value <= 4'h0; // @[Counter.scala 60:40]
    end else if (do_deq) begin // @[Decoupled.scala 233:17]
      if (wrap_1) begin // @[Counter.scala 86:20]
        deq_ptr_value <= 4'h0; // @[Counter.scala 86:28]
      end else begin
        deq_ptr_value <= _value_T_3; // @[Counter.scala 76:15]
      end
    end
    if (reset) begin // @[Decoupled.scala 221:27]
      maybe_full <= 1'h0; // @[Decoupled.scala 221:27]
    end else if (do_enq != do_deq) begin // @[Decoupled.scala 236:28]
      maybe_full <= do_enq; // @[Decoupled.scala 237:16]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_GARBAGE_ASSIGN
  _RAND_1 = {2{`RANDOM}};
  _RAND_3 = {1{`RANDOM}};
  _RAND_5 = {1{`RANDOM}};
  _RAND_7 = {1{`RANDOM}};
  _RAND_9 = {1{`RANDOM}};
  _RAND_11 = {1{`RANDOM}};
  _RAND_13 = {1{`RANDOM}};
  _RAND_15 = {1{`RANDOM}};
  _RAND_17 = {1{`RANDOM}};
  _RAND_19 = {1{`RANDOM}};
  _RAND_21 = {1{`RANDOM}};
  _RAND_23 = {1{`RANDOM}};
`endif // RANDOMIZE_GARBAGE_ASSIGN
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {2{`RANDOM}};
  for (initvar = 0; initvar < 10; initvar = initvar+1)
    ram_addr[initvar] = _RAND_0[63:0];
  _RAND_2 = {1{`RANDOM}};
  for (initvar = 0; initvar < 10; initvar = initvar+1)
    ram_len[initvar] = _RAND_2[31:0];
  _RAND_4 = {1{`RANDOM}};
  for (initvar = 0; initvar < 10; initvar = initvar+1)
    ram_eop[initvar] = _RAND_4[0:0];
  _RAND_6 = {1{`RANDOM}};
  for (initvar = 0; initvar < 10; initvar = initvar+1)
    ram_sop[initvar] = _RAND_6[0:0];
  _RAND_8 = {1{`RANDOM}};
  for (initvar = 0; initvar < 10; initvar = initvar+1)
    ram_mrkr_req[initvar] = _RAND_8[0:0];
  _RAND_10 = {1{`RANDOM}};
  for (initvar = 0; initvar < 10; initvar = initvar+1)
    ram_sdi[initvar] = _RAND_10[0:0];
  _RAND_12 = {1{`RANDOM}};
  for (initvar = 0; initvar < 10; initvar = initvar+1)
    ram_qid[initvar] = _RAND_12[10:0];
  _RAND_14 = {1{`RANDOM}};
  for (initvar = 0; initvar < 10; initvar = initvar+1)
    ram_error[initvar] = _RAND_14[0:0];
  _RAND_16 = {1{`RANDOM}};
  for (initvar = 0; initvar < 10; initvar = initvar+1)
    ram_func[initvar] = _RAND_16[7:0];
  _RAND_18 = {1{`RANDOM}};
  for (initvar = 0; initvar < 10; initvar = initvar+1)
    ram_cidx[initvar] = _RAND_18[15:0];
  _RAND_20 = {1{`RANDOM}};
  for (initvar = 0; initvar < 10; initvar = initvar+1)
    ram_port_id[initvar] = _RAND_20[2:0];
  _RAND_22 = {1{`RANDOM}};
  for (initvar = 0; initvar < 10; initvar = initvar+1)
    ram_no_dma[initvar] = _RAND_22[0:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  enq_ptr_value = _RAND_24[3:0];
  _RAND_25 = {1{`RANDOM}};
  deq_ptr_value = _RAND_25[3:0];
  _RAND_26 = {1{`RANDOM}};
  maybe_full = _RAND_26[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Queue_1(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input  [63:0] io_enq_bits_addr,
  input  [10:0] io_enq_bits_qid,
  input         io_enq_bits_error,
  input  [7:0]  io_enq_bits_func,
  input  [2:0]  io_enq_bits_port_id,
  input  [6:0]  io_enq_bits_pfch_tag,
  input  [31:0] io_enq_bits_len,
  input         io_deq_ready,
  output        io_deq_valid,
  output [63:0] io_deq_bits_addr,
  output [10:0] io_deq_bits_qid,
  output        io_deq_bits_error,
  output [7:0]  io_deq_bits_func,
  output [2:0]  io_deq_bits_port_id,
  output [6:0]  io_deq_bits_pfch_tag,
  output [31:0] io_deq_bits_len,
  output [3:0]  io_count
);
`ifdef RANDOMIZE_GARBAGE_ASSIGN
  reg [63:0] _RAND_1;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_13;
`endif // RANDOMIZE_GARBAGE_ASSIGN
`ifdef RANDOMIZE_MEM_INIT
  reg [63:0] _RAND_0;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_12;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
`endif // RANDOMIZE_REG_INIT
  reg [63:0] ram_addr [0:9]; // @[Decoupled.scala 218:16]
  wire [63:0] ram_addr_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16]
  wire [3:0] ram_addr_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16]
  wire [63:0] ram_addr_MPORT_data; // @[Decoupled.scala 218:16]
  wire [3:0] ram_addr_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_addr_MPORT_mask; // @[Decoupled.scala 218:16]
  wire  ram_addr_MPORT_en; // @[Decoupled.scala 218:16]
  reg [10:0] ram_qid [0:9]; // @[Decoupled.scala 218:16]
  wire [10:0] ram_qid_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16]
  wire [3:0] ram_qid_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16]
  wire [10:0] ram_qid_MPORT_data; // @[Decoupled.scala 218:16]
  wire [3:0] ram_qid_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_qid_MPORT_mask; // @[Decoupled.scala 218:16]
  wire  ram_qid_MPORT_en; // @[Decoupled.scala 218:16]
  reg  ram_error [0:9]; // @[Decoupled.scala 218:16]
  wire  ram_error_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16]
  wire [3:0] ram_error_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_error_MPORT_data; // @[Decoupled.scala 218:16]
  wire [3:0] ram_error_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_error_MPORT_mask; // @[Decoupled.scala 218:16]
  wire  ram_error_MPORT_en; // @[Decoupled.scala 218:16]
  reg [7:0] ram_func [0:9]; // @[Decoupled.scala 218:16]
  wire [7:0] ram_func_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16]
  wire [3:0] ram_func_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16]
  wire [7:0] ram_func_MPORT_data; // @[Decoupled.scala 218:16]
  wire [3:0] ram_func_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_func_MPORT_mask; // @[Decoupled.scala 218:16]
  wire  ram_func_MPORT_en; // @[Decoupled.scala 218:16]
  reg [2:0] ram_port_id [0:9]; // @[Decoupled.scala 218:16]
  wire [2:0] ram_port_id_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16]
  wire [3:0] ram_port_id_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16]
  wire [2:0] ram_port_id_MPORT_data; // @[Decoupled.scala 218:16]
  wire [3:0] ram_port_id_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_port_id_MPORT_mask; // @[Decoupled.scala 218:16]
  wire  ram_port_id_MPORT_en; // @[Decoupled.scala 218:16]
  reg [6:0] ram_pfch_tag [0:9]; // @[Decoupled.scala 218:16]
  wire [6:0] ram_pfch_tag_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16]
  wire [3:0] ram_pfch_tag_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16]
  wire [6:0] ram_pfch_tag_MPORT_data; // @[Decoupled.scala 218:16]
  wire [3:0] ram_pfch_tag_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_pfch_tag_MPORT_mask; // @[Decoupled.scala 218:16]
  wire  ram_pfch_tag_MPORT_en; // @[Decoupled.scala 218:16]
  reg [31:0] ram_len [0:9]; // @[Decoupled.scala 218:16]
  wire [31:0] ram_len_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16]
  wire [3:0] ram_len_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16]
  wire [31:0] ram_len_MPORT_data; // @[Decoupled.scala 218:16]
  wire [3:0] ram_len_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_len_MPORT_mask; // @[Decoupled.scala 218:16]
  wire  ram_len_MPORT_en; // @[Decoupled.scala 218:16]
  reg [3:0] enq_ptr_value; // @[Counter.scala 60:40]
  reg [3:0] deq_ptr_value; // @[Counter.scala 60:40]
  reg  maybe_full; // @[Decoupled.scala 221:27]
  wire  ptr_match = enq_ptr_value == deq_ptr_value; // @[Decoupled.scala 223:33]
  wire  empty = ptr_match & ~maybe_full; // @[Decoupled.scala 224:25]
  wire  full = ptr_match & maybe_full; // @[Decoupled.scala 225:24]
  wire  do_enq = io_enq_ready & io_enq_valid; // @[Decoupled.scala 40:37]
  wire  do_deq = io_deq_ready & io_deq_valid; // @[Decoupled.scala 40:37]
  wire  wrap = enq_ptr_value == 4'h9; // @[Counter.scala 72:24]
  wire [3:0] _value_T_1 = enq_ptr_value + 4'h1; // @[Counter.scala 76:24]
  wire  wrap_1 = deq_ptr_value == 4'h9; // @[Counter.scala 72:24]
  wire [3:0] _value_T_3 = deq_ptr_value + 4'h1; // @[Counter.scala 76:24]
  wire [3:0] ptr_diff = enq_ptr_value - deq_ptr_value; // @[Decoupled.scala 257:32]
  wire [3:0] _io_count_T = maybe_full ? 4'ha : 4'h0; // @[Decoupled.scala 262:24]
  wire [3:0] _io_count_T_3 = 4'ha + ptr_diff; // @[Decoupled.scala 265:38]
  wire [3:0] _io_count_T_4 = deq_ptr_value > enq_ptr_value ? _io_count_T_3 : ptr_diff; // @[Decoupled.scala 264:24]
  assign ram_addr_io_deq_bits_MPORT_addr = deq_ptr_value;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign ram_addr_io_deq_bits_MPORT_data = ram_addr[ram_addr_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  `else
  assign ram_addr_io_deq_bits_MPORT_data = ram_addr_io_deq_bits_MPORT_addr >= 4'ha ? _RAND_1[63:0] :
    ram_addr[ram_addr_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign ram_addr_MPORT_data = io_enq_bits_addr;
  assign ram_addr_MPORT_addr = enq_ptr_value;
  assign ram_addr_MPORT_mask = 1'h1;
  assign ram_addr_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_qid_io_deq_bits_MPORT_addr = deq_ptr_value;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign ram_qid_io_deq_bits_MPORT_data = ram_qid[ram_qid_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  `else
  assign ram_qid_io_deq_bits_MPORT_data = ram_qid_io_deq_bits_MPORT_addr >= 4'ha ? _RAND_3[10:0] :
    ram_qid[ram_qid_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign ram_qid_MPORT_data = io_enq_bits_qid;
  assign ram_qid_MPORT_addr = enq_ptr_value;
  assign ram_qid_MPORT_mask = 1'h1;
  assign ram_qid_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_error_io_deq_bits_MPORT_addr = deq_ptr_value;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign ram_error_io_deq_bits_MPORT_data = ram_error[ram_error_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  `else
  assign ram_error_io_deq_bits_MPORT_data = ram_error_io_deq_bits_MPORT_addr >= 4'ha ? _RAND_5[0:0] :
    ram_error[ram_error_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign ram_error_MPORT_data = io_enq_bits_error;
  assign ram_error_MPORT_addr = enq_ptr_value;
  assign ram_error_MPORT_mask = 1'h1;
  assign ram_error_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_func_io_deq_bits_MPORT_addr = deq_ptr_value;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign ram_func_io_deq_bits_MPORT_data = ram_func[ram_func_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  `else
  assign ram_func_io_deq_bits_MPORT_data = ram_func_io_deq_bits_MPORT_addr >= 4'ha ? _RAND_7[7:0] :
    ram_func[ram_func_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign ram_func_MPORT_data = io_enq_bits_func;
  assign ram_func_MPORT_addr = enq_ptr_value;
  assign ram_func_MPORT_mask = 1'h1;
  assign ram_func_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_port_id_io_deq_bits_MPORT_addr = deq_ptr_value;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign ram_port_id_io_deq_bits_MPORT_data = ram_port_id[ram_port_id_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  `else
  assign ram_port_id_io_deq_bits_MPORT_data = ram_port_id_io_deq_bits_MPORT_addr >= 4'ha ? _RAND_9[2:0] :
    ram_port_id[ram_port_id_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign ram_port_id_MPORT_data = io_enq_bits_port_id;
  assign ram_port_id_MPORT_addr = enq_ptr_value;
  assign ram_port_id_MPORT_mask = 1'h1;
  assign ram_port_id_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_pfch_tag_io_deq_bits_MPORT_addr = deq_ptr_value;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign ram_pfch_tag_io_deq_bits_MPORT_data = ram_pfch_tag[ram_pfch_tag_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  `else
  assign ram_pfch_tag_io_deq_bits_MPORT_data = ram_pfch_tag_io_deq_bits_MPORT_addr >= 4'ha ? _RAND_11[6:0] :
    ram_pfch_tag[ram_pfch_tag_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign ram_pfch_tag_MPORT_data = io_enq_bits_pfch_tag;
  assign ram_pfch_tag_MPORT_addr = enq_ptr_value;
  assign ram_pfch_tag_MPORT_mask = 1'h1;
  assign ram_pfch_tag_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_len_io_deq_bits_MPORT_addr = deq_ptr_value;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign ram_len_io_deq_bits_MPORT_data = ram_len[ram_len_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  `else
  assign ram_len_io_deq_bits_MPORT_data = ram_len_io_deq_bits_MPORT_addr >= 4'ha ? _RAND_13[31:0] :
    ram_len[ram_len_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign ram_len_MPORT_data = io_enq_bits_len;
  assign ram_len_MPORT_addr = enq_ptr_value;
  assign ram_len_MPORT_mask = 1'h1;
  assign ram_len_MPORT_en = io_enq_ready & io_enq_valid;
  assign io_enq_ready = ~full; // @[Decoupled.scala 241:19]
  assign io_deq_valid = ~empty; // @[Decoupled.scala 240:19]
  assign io_deq_bits_addr = ram_addr_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15]
  assign io_deq_bits_qid = ram_qid_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15]
  assign io_deq_bits_error = ram_error_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15]
  assign io_deq_bits_func = ram_func_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15]
  assign io_deq_bits_port_id = ram_port_id_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15]
  assign io_deq_bits_pfch_tag = ram_pfch_tag_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15]
  assign io_deq_bits_len = ram_len_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15]
  assign io_count = ptr_match ? _io_count_T : _io_count_T_4; // @[Decoupled.scala 261:20]
  always @(posedge clock) begin
    if(ram_addr_MPORT_en & ram_addr_MPORT_mask) begin
      ram_addr[ram_addr_MPORT_addr] <= ram_addr_MPORT_data; // @[Decoupled.scala 218:16]
    end
    if(ram_qid_MPORT_en & ram_qid_MPORT_mask) begin
      ram_qid[ram_qid_MPORT_addr] <= ram_qid_MPORT_data; // @[Decoupled.scala 218:16]
    end
    if(ram_error_MPORT_en & ram_error_MPORT_mask) begin
      ram_error[ram_error_MPORT_addr] <= ram_error_MPORT_data; // @[Decoupled.scala 218:16]
    end
    if(ram_func_MPORT_en & ram_func_MPORT_mask) begin
      ram_func[ram_func_MPORT_addr] <= ram_func_MPORT_data; // @[Decoupled.scala 218:16]
    end
    if(ram_port_id_MPORT_en & ram_port_id_MPORT_mask) begin
      ram_port_id[ram_port_id_MPORT_addr] <= ram_port_id_MPORT_data; // @[Decoupled.scala 218:16]
    end
    if(ram_pfch_tag_MPORT_en & ram_pfch_tag_MPORT_mask) begin
      ram_pfch_tag[ram_pfch_tag_MPORT_addr] <= ram_pfch_tag_MPORT_data; // @[Decoupled.scala 218:16]
    end
    if(ram_len_MPORT_en & ram_len_MPORT_mask) begin
      ram_len[ram_len_MPORT_addr] <= ram_len_MPORT_data; // @[Decoupled.scala 218:16]
    end
    if (reset) begin // @[Counter.scala 60:40]
      enq_ptr_value <= 4'h0; // @[Counter.scala 60:40]
    end else if (do_enq) begin // @[Decoupled.scala 229:17]
      if (wrap) begin // @[Counter.scala 86:20]
        enq_ptr_value <= 4'h0; // @[Counter.scala 86:28]
      end else begin
        enq_ptr_value <= _value_T_1; // @[Counter.scala 76:15]
      end
    end
    if (reset) begin // @[Counter.scala 60:40]
      deq_ptr_value <= 4'h0; // @[Counter.scala 60:40]
    end else if (do_deq) begin // @[Decoupled.scala 233:17]
      if (wrap_1) begin // @[Counter.scala 86:20]
        deq_ptr_value <= 4'h0; // @[Counter.scala 86:28]
      end else begin
        deq_ptr_value <= _value_T_3; // @[Counter.scala 76:15]
      end
    end
    if (reset) begin // @[Decoupled.scala 221:27]
      maybe_full <= 1'h0; // @[Decoupled.scala 221:27]
    end else if (do_enq != do_deq) begin // @[Decoupled.scala 236:28]
      maybe_full <= do_enq; // @[Decoupled.scala 237:16]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_GARBAGE_ASSIGN
  _RAND_1 = {2{`RANDOM}};
  _RAND_3 = {1{`RANDOM}};
  _RAND_5 = {1{`RANDOM}};
  _RAND_7 = {1{`RANDOM}};
  _RAND_9 = {1{`RANDOM}};
  _RAND_11 = {1{`RANDOM}};
  _RAND_13 = {1{`RANDOM}};
`endif // RANDOMIZE_GARBAGE_ASSIGN
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {2{`RANDOM}};
  for (initvar = 0; initvar < 10; initvar = initvar+1)
    ram_addr[initvar] = _RAND_0[63:0];
  _RAND_2 = {1{`RANDOM}};
  for (initvar = 0; initvar < 10; initvar = initvar+1)
    ram_qid[initvar] = _RAND_2[10:0];
  _RAND_4 = {1{`RANDOM}};
  for (initvar = 0; initvar < 10; initvar = initvar+1)
    ram_error[initvar] = _RAND_4[0:0];
  _RAND_6 = {1{`RANDOM}};
  for (initvar = 0; initvar < 10; initvar = initvar+1)
    ram_func[initvar] = _RAND_6[7:0];
  _RAND_8 = {1{`RANDOM}};
  for (initvar = 0; initvar < 10; initvar = initvar+1)
    ram_port_id[initvar] = _RAND_8[2:0];
  _RAND_10 = {1{`RANDOM}};
  for (initvar = 0; initvar < 10; initvar = initvar+1)
    ram_pfch_tag[initvar] = _RAND_10[6:0];
  _RAND_12 = {1{`RANDOM}};
  for (initvar = 0; initvar < 10; initvar = initvar+1)
    ram_len[initvar] = _RAND_12[31:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  enq_ptr_value = _RAND_14[3:0];
  _RAND_15 = {1{`RANDOM}};
  deq_ptr_value = _RAND_15[3:0];
  _RAND_16 = {1{`RANDOM}};
  maybe_full = _RAND_16[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module TLB(
  input         clock,
  input         reset,
  output        io__wr_tlb_ready,
  input         io__wr_tlb_valid,
  input  [31:0] io__wr_tlb_bits_vaddr_high,
  input  [31:0] io__wr_tlb_bits_vaddr_low,
  input  [31:0] io__wr_tlb_bits_paddr_high,
  input  [31:0] io__wr_tlb_bits_paddr_low,
  input         io__wr_tlb_bits_is_base,
  output        io__h2c_in_ready,
  input         io__h2c_in_valid,
  input  [63:0] io__h2c_in_bits_addr,
  input  [31:0] io__h2c_in_bits_len,
  input         io__h2c_in_bits_eop,
  input         io__h2c_in_bits_sop,
  input         io__h2c_in_bits_mrkr_req,
  input         io__h2c_in_bits_sdi,
  input  [10:0] io__h2c_in_bits_qid,
  input         io__h2c_in_bits_error,
  input  [7:0]  io__h2c_in_bits_func,
  input  [15:0] io__h2c_in_bits_cidx,
  input  [2:0]  io__h2c_in_bits_port_id,
  input         io__h2c_in_bits_no_dma,
  output        io__c2h_in_ready,
  input         io__c2h_in_valid,
  input  [63:0] io__c2h_in_bits_addr,
  input  [10:0] io__c2h_in_bits_qid,
  input         io__c2h_in_bits_error,
  input  [7:0]  io__c2h_in_bits_func,
  input  [2:0]  io__c2h_in_bits_port_id,
  input  [6:0]  io__c2h_in_bits_pfch_tag,
  input  [31:0] io__c2h_in_bits_len,
  input         io__h2c_out_ready,
  output        io__h2c_out_valid,
  output [63:0] io__h2c_out_bits_addr,
  output [31:0] io__h2c_out_bits_len,
  output        io__h2c_out_bits_eop,
  output        io__h2c_out_bits_sop,
  output        io__h2c_out_bits_mrkr_req,
  output        io__h2c_out_bits_sdi,
  output [10:0] io__h2c_out_bits_qid,
  output        io__h2c_out_bits_error,
  output [7:0]  io__h2c_out_bits_func,
  output [15:0] io__h2c_out_bits_cidx,
  output [2:0]  io__h2c_out_bits_port_id,
  output        io__h2c_out_bits_no_dma,
  input         io__c2h_out_ready,
  output        io__c2h_out_valid,
  output [63:0] io__c2h_out_bits_addr,
  output [10:0] io__c2h_out_bits_qid,
  output        io__c2h_out_bits_error,
  output [7:0]  io__c2h_out_bits_func,
  output [2:0]  io__c2h_out_bits_port_id,
  output [6:0]  io__c2h_out_bits_pfch_tag,
  output [31:0] io__c2h_out_bits_len,
  output [31:0] io__tlb_miss_count,
  output [31:0] io_tlb_miss_count
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
`endif // RANDOMIZE_REG_INIT
  wire  tlb_table_clock; // @[XRam.scala 102:23]
  wire  tlb_table_reset; // @[XRam.scala 102:23]
  wire [12:0] tlb_table_io_addr_a; // @[XRam.scala 102:23]
  wire [12:0] tlb_table_io_addr_b; // @[XRam.scala 102:23]
  wire  tlb_table_io_wr_en_a; // @[XRam.scala 102:23]
  wire [63:0] tlb_table_io_data_in_a; // @[XRam.scala 102:23]
  wire [63:0] tlb_table_io_data_out_a; // @[XRam.scala 102:23]
  wire [63:0] tlb_table_io_data_out_b; // @[XRam.scala 102:23]
  wire  q_h2c_clock; // @[TLB.scala 74:57]
  wire  q_h2c_reset; // @[TLB.scala 74:57]
  wire  q_h2c_io_enq_ready; // @[TLB.scala 74:57]
  wire  q_h2c_io_enq_valid; // @[TLB.scala 74:57]
  wire [63:0] q_h2c_io_enq_bits_addr; // @[TLB.scala 74:57]
  wire [31:0] q_h2c_io_enq_bits_len; // @[TLB.scala 74:57]
  wire  q_h2c_io_enq_bits_eop; // @[TLB.scala 74:57]
  wire  q_h2c_io_enq_bits_sop; // @[TLB.scala 74:57]
  wire  q_h2c_io_enq_bits_mrkr_req; // @[TLB.scala 74:57]
  wire  q_h2c_io_enq_bits_sdi; // @[TLB.scala 74:57]
  wire [10:0] q_h2c_io_enq_bits_qid; // @[TLB.scala 74:57]
  wire  q_h2c_io_enq_bits_error; // @[TLB.scala 74:57]
  wire [7:0] q_h2c_io_enq_bits_func; // @[TLB.scala 74:57]
  wire [15:0] q_h2c_io_enq_bits_cidx; // @[TLB.scala 74:57]
  wire [2:0] q_h2c_io_enq_bits_port_id; // @[TLB.scala 74:57]
  wire  q_h2c_io_enq_bits_no_dma; // @[TLB.scala 74:57]
  wire  q_h2c_io_deq_ready; // @[TLB.scala 74:57]
  wire  q_h2c_io_deq_valid; // @[TLB.scala 74:57]
  wire [63:0] q_h2c_io_deq_bits_addr; // @[TLB.scala 74:57]
  wire [31:0] q_h2c_io_deq_bits_len; // @[TLB.scala 74:57]
  wire  q_h2c_io_deq_bits_eop; // @[TLB.scala 74:57]
  wire  q_h2c_io_deq_bits_sop; // @[TLB.scala 74:57]
  wire  q_h2c_io_deq_bits_mrkr_req; // @[TLB.scala 74:57]
  wire  q_h2c_io_deq_bits_sdi; // @[TLB.scala 74:57]
  wire [10:0] q_h2c_io_deq_bits_qid; // @[TLB.scala 74:57]
  wire  q_h2c_io_deq_bits_error; // @[TLB.scala 74:57]
  wire [7:0] q_h2c_io_deq_bits_func; // @[TLB.scala 74:57]
  wire [15:0] q_h2c_io_deq_bits_cidx; // @[TLB.scala 74:57]
  wire [2:0] q_h2c_io_deq_bits_port_id; // @[TLB.scala 74:57]
  wire  q_h2c_io_deq_bits_no_dma; // @[TLB.scala 74:57]
  wire [3:0] q_h2c_io_count; // @[TLB.scala 74:57]
  wire  q_c2h_clock; // @[TLB.scala 75:57]
  wire  q_c2h_reset; // @[TLB.scala 75:57]
  wire  q_c2h_io_enq_ready; // @[TLB.scala 75:57]
  wire  q_c2h_io_enq_valid; // @[TLB.scala 75:57]
  wire [63:0] q_c2h_io_enq_bits_addr; // @[TLB.scala 75:57]
  wire [10:0] q_c2h_io_enq_bits_qid; // @[TLB.scala 75:57]
  wire  q_c2h_io_enq_bits_error; // @[TLB.scala 75:57]
  wire [7:0] q_c2h_io_enq_bits_func; // @[TLB.scala 75:57]
  wire [2:0] q_c2h_io_enq_bits_port_id; // @[TLB.scala 75:57]
  wire [6:0] q_c2h_io_enq_bits_pfch_tag; // @[TLB.scala 75:57]
  wire [31:0] q_c2h_io_enq_bits_len; // @[TLB.scala 75:57]
  wire  q_c2h_io_deq_ready; // @[TLB.scala 75:57]
  wire  q_c2h_io_deq_valid; // @[TLB.scala 75:57]
  wire [63:0] q_c2h_io_deq_bits_addr; // @[TLB.scala 75:57]
  wire [10:0] q_c2h_io_deq_bits_qid; // @[TLB.scala 75:57]
  wire  q_c2h_io_deq_bits_error; // @[TLB.scala 75:57]
  wire [7:0] q_c2h_io_deq_bits_func; // @[TLB.scala 75:57]
  wire [2:0] q_c2h_io_deq_bits_port_id; // @[TLB.scala 75:57]
  wire [6:0] q_c2h_io_deq_bits_pfch_tag; // @[TLB.scala 75:57]
  wire [31:0] q_c2h_io_deq_bits_len; // @[TLB.scala 75:57]
  wire [3:0] q_c2h_io_count; // @[TLB.scala 75:57]
  reg [42:0] base_page; // @[TLB.scala 37:50]
  reg [31:0] tlb_miss_count; // @[TLB.scala 38:50]
  reg [13:0] wrtlb_index; // @[TLB.scala 40:50]
  wire [42:0] h2c_page = io__h2c_in_bits_addr[63:21]; // @[TLB.scala 41:62]
  wire [42:0] h2c_index = h2c_page - base_page; // @[TLB.scala 42:52]
  wire [42:0] _GEN_12 = {{29'd0}, wrtlb_index}; // @[TLB.scala 43:90]
  wire [42:0] _h2c_outrange_T_2 = base_page + _GEN_12; // @[TLB.scala 43:90]
  wire  h2c_outrange = h2c_page < base_page | h2c_page >= _h2c_outrange_T_2; // @[TLB.scala 43:66]
  wire [42:0] c2h_page = io__c2h_in_bits_addr[63:21]; // @[TLB.scala 44:62]
  wire [42:0] c2h_index = c2h_page - base_page; // @[TLB.scala 45:52]
  wire  c2h_outrange = c2h_page < base_page | c2h_page >= _h2c_outrange_T_2; // @[TLB.scala 46:66]
  wire  _tlb_table_io_wr_en_a_T = io__wr_tlb_ready & io__wr_tlb_valid; // @[Decoupled.scala 40:37]
  wire [13:0] _wrtlb_index_T_1 = wrtlb_index + 14'h1; // @[TLB.scala 56:72]
  wire [63:0] _base_page_T = {io__wr_tlb_bits_vaddr_high,io__wr_tlb_bits_vaddr_low}; // @[Cat.scala 30:58]
  wire [13:0] _GEN_1 = io__wr_tlb_bits_is_base ? 14'h0 : wrtlb_index; // @[TLB.scala 57:51 TLB.scala 59:49 TLB.scala 55:49]
  wire [42:0] _GEN_4 = _tlb_table_io_wr_en_a_T ? {{29'd0}, _GEN_1} : h2c_index; // @[TLB.scala 54:31 TLB.scala 64:41]
  reg [31:0] h2c_bits_delay_REG_len; // @[TLB.scala 70:59]
  reg  h2c_bits_delay_REG_eop; // @[TLB.scala 70:59]
  reg  h2c_bits_delay_REG_sop; // @[TLB.scala 70:59]
  reg  h2c_bits_delay_REG_mrkr_req; // @[TLB.scala 70:59]
  reg  h2c_bits_delay_REG_sdi; // @[TLB.scala 70:59]
  reg [10:0] h2c_bits_delay_REG_qid; // @[TLB.scala 70:59]
  reg  h2c_bits_delay_REG_error; // @[TLB.scala 70:59]
  reg [7:0] h2c_bits_delay_REG_func; // @[TLB.scala 70:59]
  reg [15:0] h2c_bits_delay_REG_cidx; // @[TLB.scala 70:59]
  reg [2:0] h2c_bits_delay_REG_port_id; // @[TLB.scala 70:59]
  reg  h2c_bits_delay_REG_no_dma; // @[TLB.scala 70:59]
  reg [31:0] h2c_bits_delay_REG_1_len; // @[TLB.scala 70:51]
  reg  h2c_bits_delay_REG_1_eop; // @[TLB.scala 70:51]
  reg  h2c_bits_delay_REG_1_sop; // @[TLB.scala 70:51]
  reg  h2c_bits_delay_REG_1_mrkr_req; // @[TLB.scala 70:51]
  reg  h2c_bits_delay_REG_1_sdi; // @[TLB.scala 70:51]
  reg [10:0] h2c_bits_delay_REG_1_qid; // @[TLB.scala 70:51]
  reg  h2c_bits_delay_REG_1_error; // @[TLB.scala 70:51]
  reg [7:0] h2c_bits_delay_REG_1_func; // @[TLB.scala 70:51]
  reg [15:0] h2c_bits_delay_REG_1_cidx; // @[TLB.scala 70:51]
  reg [2:0] h2c_bits_delay_REG_1_port_id; // @[TLB.scala 70:51]
  reg  h2c_bits_delay_REG_1_no_dma; // @[TLB.scala 70:51]
  reg [10:0] c2h_bits_delay_REG_qid; // @[TLB.scala 71:59]
  reg  c2h_bits_delay_REG_error; // @[TLB.scala 71:59]
  reg [7:0] c2h_bits_delay_REG_func; // @[TLB.scala 71:59]
  reg [2:0] c2h_bits_delay_REG_port_id; // @[TLB.scala 71:59]
  reg [6:0] c2h_bits_delay_REG_pfch_tag; // @[TLB.scala 71:59]
  reg [31:0] c2h_bits_delay_REG_len; // @[TLB.scala 71:59]
  reg [10:0] c2h_bits_delay_REG_1_qid; // @[TLB.scala 71:51]
  reg  c2h_bits_delay_REG_1_error; // @[TLB.scala 71:51]
  reg [7:0] c2h_bits_delay_REG_1_func; // @[TLB.scala 71:51]
  reg [2:0] c2h_bits_delay_REG_1_port_id; // @[TLB.scala 71:51]
  reg [6:0] c2h_bits_delay_REG_1_pfch_tag; // @[TLB.scala 71:51]
  reg [31:0] c2h_bits_delay_REG_1_len; // @[TLB.scala 71:51]
  reg [20:0] h2c_bits_delay_addr_REG; // @[TLB.scala 72:77]
  reg [20:0] h2c_bits_delay_addr_REG_1; // @[TLB.scala 72:69]
  wire [63:0] _GEN_14 = {{43'd0}, h2c_bits_delay_addr_REG_1}; // @[TLB.scala 72:60]
  reg [20:0] c2h_bits_delay_addr_REG; // @[TLB.scala 73:77]
  reg [20:0] c2h_bits_delay_addr_REG_1; // @[TLB.scala 73:69]
  wire [63:0] _GEN_15 = {{43'd0}, c2h_bits_delay_addr_REG_1}; // @[TLB.scala 73:60]
  reg  REG; // @[TLB.scala 80:29]
  reg  REG_1; // @[TLB.scala 80:21]
  reg  REG_2; // @[TLB.scala 80:66]
  reg  REG_3; // @[TLB.scala 80:58]
  reg  REG_4; // @[TLB.scala 80:104]
  reg  REG_5; // @[TLB.scala 80:96]
  reg  REG_6; // @[TLB.scala 86:29]
  reg  REG_7; // @[TLB.scala 86:21]
  reg  REG_8; // @[TLB.scala 86:66]
  reg  REG_9; // @[TLB.scala 86:58]
  reg  REG_10; // @[TLB.scala 86:104]
  reg  REG_11; // @[TLB.scala 86:96]
  wire  h2c_miss = h2c_outrange & io__h2c_in_valid & io__h2c_in_ready; // @[TLB.scala 92:58]
  wire  c2h_miss = c2h_outrange & io__c2h_in_valid & io__c2h_in_ready; // @[TLB.scala 93:58]
  wire [31:0] _tlb_miss_count_T_1 = tlb_miss_count + 32'h1; // @[TLB.scala 95:50]
  wire [31:0] _tlb_miss_count_T_3 = tlb_miss_count + 32'h2; // @[TLB.scala 97:58]
  XRam tlb_table ( // @[XRam.scala 102:23]
    .clock(tlb_table_clock),
    .reset(tlb_table_reset),
    .io_addr_a(tlb_table_io_addr_a),
    .io_addr_b(tlb_table_io_addr_b),
    .io_wr_en_a(tlb_table_io_wr_en_a),
    .io_data_in_a(tlb_table_io_data_in_a),
    .io_data_out_a(tlb_table_io_data_out_a),
    .io_data_out_b(tlb_table_io_data_out_b)
  );
  Queue q_h2c ( // @[TLB.scala 74:57]
    .clock(q_h2c_clock),
    .reset(q_h2c_reset),
    .io_enq_ready(q_h2c_io_enq_ready),
    .io_enq_valid(q_h2c_io_enq_valid),
    .io_enq_bits_addr(q_h2c_io_enq_bits_addr),
    .io_enq_bits_len(q_h2c_io_enq_bits_len),
    .io_enq_bits_eop(q_h2c_io_enq_bits_eop),
    .io_enq_bits_sop(q_h2c_io_enq_bits_sop),
    .io_enq_bits_mrkr_req(q_h2c_io_enq_bits_mrkr_req),
    .io_enq_bits_sdi(q_h2c_io_enq_bits_sdi),
    .io_enq_bits_qid(q_h2c_io_enq_bits_qid),
    .io_enq_bits_error(q_h2c_io_enq_bits_error),
    .io_enq_bits_func(q_h2c_io_enq_bits_func),
    .io_enq_bits_cidx(q_h2c_io_enq_bits_cidx),
    .io_enq_bits_port_id(q_h2c_io_enq_bits_port_id),
    .io_enq_bits_no_dma(q_h2c_io_enq_bits_no_dma),
    .io_deq_ready(q_h2c_io_deq_ready),
    .io_deq_valid(q_h2c_io_deq_valid),
    .io_deq_bits_addr(q_h2c_io_deq_bits_addr),
    .io_deq_bits_len(q_h2c_io_deq_bits_len),
    .io_deq_bits_eop(q_h2c_io_deq_bits_eop),
    .io_deq_bits_sop(q_h2c_io_deq_bits_sop),
    .io_deq_bits_mrkr_req(q_h2c_io_deq_bits_mrkr_req),
    .io_deq_bits_sdi(q_h2c_io_deq_bits_sdi),
    .io_deq_bits_qid(q_h2c_io_deq_bits_qid),
    .io_deq_bits_error(q_h2c_io_deq_bits_error),
    .io_deq_bits_func(q_h2c_io_deq_bits_func),
    .io_deq_bits_cidx(q_h2c_io_deq_bits_cidx),
    .io_deq_bits_port_id(q_h2c_io_deq_bits_port_id),
    .io_deq_bits_no_dma(q_h2c_io_deq_bits_no_dma),
    .io_count(q_h2c_io_count)
  );
  Queue_1 q_c2h ( // @[TLB.scala 75:57]
    .clock(q_c2h_clock),
    .reset(q_c2h_reset),
    .io_enq_ready(q_c2h_io_enq_ready),
    .io_enq_valid(q_c2h_io_enq_valid),
    .io_enq_bits_addr(q_c2h_io_enq_bits_addr),
    .io_enq_bits_qid(q_c2h_io_enq_bits_qid),
    .io_enq_bits_error(q_c2h_io_enq_bits_error),
    .io_enq_bits_func(q_c2h_io_enq_bits_func),
    .io_enq_bits_port_id(q_c2h_io_enq_bits_port_id),
    .io_enq_bits_pfch_tag(q_c2h_io_enq_bits_pfch_tag),
    .io_enq_bits_len(q_c2h_io_enq_bits_len),
    .io_deq_ready(q_c2h_io_deq_ready),
    .io_deq_valid(q_c2h_io_deq_valid),
    .io_deq_bits_addr(q_c2h_io_deq_bits_addr),
    .io_deq_bits_qid(q_c2h_io_deq_bits_qid),
    .io_deq_bits_error(q_c2h_io_deq_bits_error),
    .io_deq_bits_func(q_c2h_io_deq_bits_func),
    .io_deq_bits_port_id(q_c2h_io_deq_bits_port_id),
    .io_deq_bits_pfch_tag(q_c2h_io_deq_bits_pfch_tag),
    .io_deq_bits_len(q_c2h_io_deq_bits_len),
    .io_count(q_c2h_io_count)
  );
  assign io__wr_tlb_ready = 1'h1; // @[TLB.scala 50:41]
  assign io__h2c_in_ready = q_h2c_io_count < 4'h8; // @[TLB.scala 77:58]
  assign io__c2h_in_ready = q_c2h_io_count < 4'h8; // @[TLB.scala 78:59]
  assign io__h2c_out_valid = q_h2c_io_deq_valid; // @[TLB.scala 102:41]
  assign io__h2c_out_bits_addr = q_h2c_io_deq_bits_addr; // @[TLB.scala 102:41]
  assign io__h2c_out_bits_len = q_h2c_io_deq_bits_len; // @[TLB.scala 102:41]
  assign io__h2c_out_bits_eop = q_h2c_io_deq_bits_eop; // @[TLB.scala 102:41]
  assign io__h2c_out_bits_sop = q_h2c_io_deq_bits_sop; // @[TLB.scala 102:41]
  assign io__h2c_out_bits_mrkr_req = q_h2c_io_deq_bits_mrkr_req; // @[TLB.scala 102:41]
  assign io__h2c_out_bits_sdi = q_h2c_io_deq_bits_sdi; // @[TLB.scala 102:41]
  assign io__h2c_out_bits_qid = q_h2c_io_deq_bits_qid; // @[TLB.scala 102:41]
  assign io__h2c_out_bits_error = q_h2c_io_deq_bits_error; // @[TLB.scala 102:41]
  assign io__h2c_out_bits_func = q_h2c_io_deq_bits_func; // @[TLB.scala 102:41]
  assign io__h2c_out_bits_cidx = q_h2c_io_deq_bits_cidx; // @[TLB.scala 102:41]
  assign io__h2c_out_bits_port_id = q_h2c_io_deq_bits_port_id; // @[TLB.scala 102:41]
  assign io__h2c_out_bits_no_dma = q_h2c_io_deq_bits_no_dma; // @[TLB.scala 102:41]
  assign io__c2h_out_valid = q_c2h_io_deq_valid; // @[TLB.scala 105:41]
  assign io__c2h_out_bits_addr = q_c2h_io_deq_bits_addr; // @[TLB.scala 105:41]
  assign io__c2h_out_bits_qid = q_c2h_io_deq_bits_qid; // @[TLB.scala 105:41]
  assign io__c2h_out_bits_error = q_c2h_io_deq_bits_error; // @[TLB.scala 105:41]
  assign io__c2h_out_bits_func = q_c2h_io_deq_bits_func; // @[TLB.scala 105:41]
  assign io__c2h_out_bits_port_id = q_c2h_io_deq_bits_port_id; // @[TLB.scala 105:41]
  assign io__c2h_out_bits_pfch_tag = q_c2h_io_deq_bits_pfch_tag; // @[TLB.scala 105:41]
  assign io__c2h_out_bits_len = q_c2h_io_deq_bits_len; // @[TLB.scala 105:41]
  assign io__tlb_miss_count = tlb_miss_count; // @[TLB.scala 107:33]
  assign io_tlb_miss_count = io__tlb_miss_count;
  assign tlb_table_clock = clock;
  assign tlb_table_reset = reset;
  assign tlb_table_io_addr_a = _GEN_4[12:0];
  assign tlb_table_io_addr_b = c2h_index[12:0]; // @[TLB.scala 66:41]
  assign tlb_table_io_wr_en_a = io__wr_tlb_ready & io__wr_tlb_valid; // @[Decoupled.scala 40:37]
  assign tlb_table_io_data_in_a = {io__wr_tlb_bits_paddr_high,io__wr_tlb_bits_paddr_low}; // @[Cat.scala 30:58]
  assign q_h2c_clock = clock;
  assign q_h2c_reset = reset;
  assign q_h2c_io_enq_valid = REG_1 & REG_3 & ~REG_5; // @[TLB.scala 80:85]
  assign q_h2c_io_enq_bits_addr = tlb_table_io_data_out_a + _GEN_14; // @[TLB.scala 72:60]
  assign q_h2c_io_enq_bits_len = h2c_bits_delay_REG_1_len; // @[TLB.scala 68:47 TLB.scala 70:41]
  assign q_h2c_io_enq_bits_eop = h2c_bits_delay_REG_1_eop; // @[TLB.scala 68:47 TLB.scala 70:41]
  assign q_h2c_io_enq_bits_sop = h2c_bits_delay_REG_1_sop; // @[TLB.scala 68:47 TLB.scala 70:41]
  assign q_h2c_io_enq_bits_mrkr_req = h2c_bits_delay_REG_1_mrkr_req; // @[TLB.scala 68:47 TLB.scala 70:41]
  assign q_h2c_io_enq_bits_sdi = h2c_bits_delay_REG_1_sdi; // @[TLB.scala 68:47 TLB.scala 70:41]
  assign q_h2c_io_enq_bits_qid = h2c_bits_delay_REG_1_qid; // @[TLB.scala 68:47 TLB.scala 70:41]
  assign q_h2c_io_enq_bits_error = h2c_bits_delay_REG_1_error; // @[TLB.scala 68:47 TLB.scala 70:41]
  assign q_h2c_io_enq_bits_func = h2c_bits_delay_REG_1_func; // @[TLB.scala 68:47 TLB.scala 70:41]
  assign q_h2c_io_enq_bits_cidx = h2c_bits_delay_REG_1_cidx; // @[TLB.scala 68:47 TLB.scala 70:41]
  assign q_h2c_io_enq_bits_port_id = h2c_bits_delay_REG_1_port_id; // @[TLB.scala 68:47 TLB.scala 70:41]
  assign q_h2c_io_enq_bits_no_dma = h2c_bits_delay_REG_1_no_dma; // @[TLB.scala 68:47 TLB.scala 70:41]
  assign q_h2c_io_deq_ready = io__h2c_out_ready; // @[TLB.scala 102:41]
  assign q_c2h_clock = clock;
  assign q_c2h_reset = reset;
  assign q_c2h_io_enq_valid = REG_7 & REG_9 & ~REG_11; // @[TLB.scala 86:85]
  assign q_c2h_io_enq_bits_addr = tlb_table_io_data_out_b + _GEN_15; // @[TLB.scala 73:60]
  assign q_c2h_io_enq_bits_qid = c2h_bits_delay_REG_1_qid; // @[TLB.scala 69:47 TLB.scala 71:41]
  assign q_c2h_io_enq_bits_error = c2h_bits_delay_REG_1_error; // @[TLB.scala 69:47 TLB.scala 71:41]
  assign q_c2h_io_enq_bits_func = c2h_bits_delay_REG_1_func; // @[TLB.scala 69:47 TLB.scala 71:41]
  assign q_c2h_io_enq_bits_port_id = c2h_bits_delay_REG_1_port_id; // @[TLB.scala 69:47 TLB.scala 71:41]
  assign q_c2h_io_enq_bits_pfch_tag = c2h_bits_delay_REG_1_pfch_tag; // @[TLB.scala 69:47 TLB.scala 71:41]
  assign q_c2h_io_enq_bits_len = c2h_bits_delay_REG_1_len; // @[TLB.scala 69:47 TLB.scala 71:41]
  assign q_c2h_io_deq_ready = io__c2h_out_ready; // @[TLB.scala 105:41]
  always @(posedge clock) begin
    if (reset) begin // @[TLB.scala 37:50]
      base_page <= 43'h0; // @[TLB.scala 37:50]
    end else if (_tlb_table_io_wr_en_a_T) begin // @[TLB.scala 54:31]
      if (io__wr_tlb_bits_is_base) begin // @[TLB.scala 57:51]
        base_page <= _base_page_T[63:21]; // @[TLB.scala 58:57]
      end
    end
    if (reset) begin // @[TLB.scala 38:50]
      tlb_miss_count <= 32'h0; // @[TLB.scala 38:50]
    end else if (h2c_miss | c2h_miss) begin // @[TLB.scala 94:34]
      if (h2c_miss & c2h_miss) begin // @[TLB.scala 96:42]
        tlb_miss_count <= _tlb_miss_count_T_3; // @[TLB.scala 97:41]
      end else begin
        tlb_miss_count <= _tlb_miss_count_T_1; // @[TLB.scala 95:33]
      end
    end else if (_tlb_table_io_wr_en_a_T) begin // @[TLB.scala 54:31]
      if (io__wr_tlb_bits_is_base) begin // @[TLB.scala 57:51]
        tlb_miss_count <= 32'h0; // @[TLB.scala 61:49]
      end
    end
    if (reset) begin // @[TLB.scala 40:50]
      wrtlb_index <= 14'h0; // @[TLB.scala 40:50]
    end else if (_tlb_table_io_wr_en_a_T) begin // @[TLB.scala 54:31]
      if (io__wr_tlb_bits_is_base) begin // @[TLB.scala 57:51]
        wrtlb_index <= 14'h1; // @[TLB.scala 60:57]
      end else begin
        wrtlb_index <= _wrtlb_index_T_1; // @[TLB.scala 56:57]
      end
    end
    h2c_bits_delay_REG_len <= io__h2c_in_bits_len; // @[TLB.scala 70:59]
    h2c_bits_delay_REG_eop <= io__h2c_in_bits_eop; // @[TLB.scala 70:59]
    h2c_bits_delay_REG_sop <= io__h2c_in_bits_sop; // @[TLB.scala 70:59]
    h2c_bits_delay_REG_mrkr_req <= io__h2c_in_bits_mrkr_req; // @[TLB.scala 70:59]
    h2c_bits_delay_REG_sdi <= io__h2c_in_bits_sdi; // @[TLB.scala 70:59]
    h2c_bits_delay_REG_qid <= io__h2c_in_bits_qid; // @[TLB.scala 70:59]
    h2c_bits_delay_REG_error <= io__h2c_in_bits_error; // @[TLB.scala 70:59]
    h2c_bits_delay_REG_func <= io__h2c_in_bits_func; // @[TLB.scala 70:59]
    h2c_bits_delay_REG_cidx <= io__h2c_in_bits_cidx; // @[TLB.scala 70:59]
    h2c_bits_delay_REG_port_id <= io__h2c_in_bits_port_id; // @[TLB.scala 70:59]
    h2c_bits_delay_REG_no_dma <= io__h2c_in_bits_no_dma; // @[TLB.scala 70:59]
    h2c_bits_delay_REG_1_len <= h2c_bits_delay_REG_len; // @[TLB.scala 70:51]
    h2c_bits_delay_REG_1_eop <= h2c_bits_delay_REG_eop; // @[TLB.scala 70:51]
    h2c_bits_delay_REG_1_sop <= h2c_bits_delay_REG_sop; // @[TLB.scala 70:51]
    h2c_bits_delay_REG_1_mrkr_req <= h2c_bits_delay_REG_mrkr_req; // @[TLB.scala 70:51]
    h2c_bits_delay_REG_1_sdi <= h2c_bits_delay_REG_sdi; // @[TLB.scala 70:51]
    h2c_bits_delay_REG_1_qid <= h2c_bits_delay_REG_qid; // @[TLB.scala 70:51]
    h2c_bits_delay_REG_1_error <= h2c_bits_delay_REG_error; // @[TLB.scala 70:51]
    h2c_bits_delay_REG_1_func <= h2c_bits_delay_REG_func; // @[TLB.scala 70:51]
    h2c_bits_delay_REG_1_cidx <= h2c_bits_delay_REG_cidx; // @[TLB.scala 70:51]
    h2c_bits_delay_REG_1_port_id <= h2c_bits_delay_REG_port_id; // @[TLB.scala 70:51]
    h2c_bits_delay_REG_1_no_dma <= h2c_bits_delay_REG_no_dma; // @[TLB.scala 70:51]
    c2h_bits_delay_REG_qid <= io__c2h_in_bits_qid; // @[TLB.scala 71:59]
    c2h_bits_delay_REG_error <= io__c2h_in_bits_error; // @[TLB.scala 71:59]
    c2h_bits_delay_REG_func <= io__c2h_in_bits_func; // @[TLB.scala 71:59]
    c2h_bits_delay_REG_port_id <= io__c2h_in_bits_port_id; // @[TLB.scala 71:59]
    c2h_bits_delay_REG_pfch_tag <= io__c2h_in_bits_pfch_tag; // @[TLB.scala 71:59]
    c2h_bits_delay_REG_len <= io__c2h_in_bits_len; // @[TLB.scala 71:59]
    c2h_bits_delay_REG_1_qid <= c2h_bits_delay_REG_qid; // @[TLB.scala 71:51]
    c2h_bits_delay_REG_1_error <= c2h_bits_delay_REG_error; // @[TLB.scala 71:51]
    c2h_bits_delay_REG_1_func <= c2h_bits_delay_REG_func; // @[TLB.scala 71:51]
    c2h_bits_delay_REG_1_port_id <= c2h_bits_delay_REG_port_id; // @[TLB.scala 71:51]
    c2h_bits_delay_REG_1_pfch_tag <= c2h_bits_delay_REG_pfch_tag; // @[TLB.scala 71:51]
    c2h_bits_delay_REG_1_len <= c2h_bits_delay_REG_len; // @[TLB.scala 71:51]
    h2c_bits_delay_addr_REG <= io__h2c_in_bits_addr[20:0]; // @[TLB.scala 72:97]
    h2c_bits_delay_addr_REG_1 <= h2c_bits_delay_addr_REG; // @[TLB.scala 72:69]
    c2h_bits_delay_addr_REG <= io__c2h_in_bits_addr[20:0]; // @[TLB.scala 73:97]
    c2h_bits_delay_addr_REG_1 <= c2h_bits_delay_addr_REG; // @[TLB.scala 73:69]
    REG <= io__h2c_in_valid; // @[TLB.scala 80:29]
    REG_1 <= REG; // @[TLB.scala 80:21]
    REG_2 <= io__h2c_in_ready; // @[TLB.scala 80:66]
    REG_3 <= REG_2; // @[TLB.scala 80:58]
    REG_4 <= h2c_page < base_page | h2c_page >= _h2c_outrange_T_2; // @[TLB.scala 43:66]
    REG_5 <= REG_4; // @[TLB.scala 80:96]
    REG_6 <= io__c2h_in_valid; // @[TLB.scala 86:29]
    REG_7 <= REG_6; // @[TLB.scala 86:21]
    REG_8 <= io__c2h_in_ready; // @[TLB.scala 86:66]
    REG_9 <= REG_8; // @[TLB.scala 86:58]
    REG_10 <= c2h_page < base_page | c2h_page >= _h2c_outrange_T_2; // @[TLB.scala 46:66]
    REG_11 <= REG_10; // @[TLB.scala 86:96]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  base_page = _RAND_0[42:0];
  _RAND_1 = {1{`RANDOM}};
  tlb_miss_count = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  wrtlb_index = _RAND_2[13:0];
  _RAND_3 = {1{`RANDOM}};
  h2c_bits_delay_REG_len = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  h2c_bits_delay_REG_eop = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  h2c_bits_delay_REG_sop = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  h2c_bits_delay_REG_mrkr_req = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  h2c_bits_delay_REG_sdi = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  h2c_bits_delay_REG_qid = _RAND_8[10:0];
  _RAND_9 = {1{`RANDOM}};
  h2c_bits_delay_REG_error = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  h2c_bits_delay_REG_func = _RAND_10[7:0];
  _RAND_11 = {1{`RANDOM}};
  h2c_bits_delay_REG_cidx = _RAND_11[15:0];
  _RAND_12 = {1{`RANDOM}};
  h2c_bits_delay_REG_port_id = _RAND_12[2:0];
  _RAND_13 = {1{`RANDOM}};
  h2c_bits_delay_REG_no_dma = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  h2c_bits_delay_REG_1_len = _RAND_14[31:0];
  _RAND_15 = {1{`RANDOM}};
  h2c_bits_delay_REG_1_eop = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  h2c_bits_delay_REG_1_sop = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  h2c_bits_delay_REG_1_mrkr_req = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  h2c_bits_delay_REG_1_sdi = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  h2c_bits_delay_REG_1_qid = _RAND_19[10:0];
  _RAND_20 = {1{`RANDOM}};
  h2c_bits_delay_REG_1_error = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  h2c_bits_delay_REG_1_func = _RAND_21[7:0];
  _RAND_22 = {1{`RANDOM}};
  h2c_bits_delay_REG_1_cidx = _RAND_22[15:0];
  _RAND_23 = {1{`RANDOM}};
  h2c_bits_delay_REG_1_port_id = _RAND_23[2:0];
  _RAND_24 = {1{`RANDOM}};
  h2c_bits_delay_REG_1_no_dma = _RAND_24[0:0];
  _RAND_25 = {1{`RANDOM}};
  c2h_bits_delay_REG_qid = _RAND_25[10:0];
  _RAND_26 = {1{`RANDOM}};
  c2h_bits_delay_REG_error = _RAND_26[0:0];
  _RAND_27 = {1{`RANDOM}};
  c2h_bits_delay_REG_func = _RAND_27[7:0];
  _RAND_28 = {1{`RANDOM}};
  c2h_bits_delay_REG_port_id = _RAND_28[2:0];
  _RAND_29 = {1{`RANDOM}};
  c2h_bits_delay_REG_pfch_tag = _RAND_29[6:0];
  _RAND_30 = {1{`RANDOM}};
  c2h_bits_delay_REG_len = _RAND_30[31:0];
  _RAND_31 = {1{`RANDOM}};
  c2h_bits_delay_REG_1_qid = _RAND_31[10:0];
  _RAND_32 = {1{`RANDOM}};
  c2h_bits_delay_REG_1_error = _RAND_32[0:0];
  _RAND_33 = {1{`RANDOM}};
  c2h_bits_delay_REG_1_func = _RAND_33[7:0];
  _RAND_34 = {1{`RANDOM}};
  c2h_bits_delay_REG_1_port_id = _RAND_34[2:0];
  _RAND_35 = {1{`RANDOM}};
  c2h_bits_delay_REG_1_pfch_tag = _RAND_35[6:0];
  _RAND_36 = {1{`RANDOM}};
  c2h_bits_delay_REG_1_len = _RAND_36[31:0];
  _RAND_37 = {1{`RANDOM}};
  h2c_bits_delay_addr_REG = _RAND_37[20:0];
  _RAND_38 = {1{`RANDOM}};
  h2c_bits_delay_addr_REG_1 = _RAND_38[20:0];
  _RAND_39 = {1{`RANDOM}};
  c2h_bits_delay_addr_REG = _RAND_39[20:0];
  _RAND_40 = {1{`RANDOM}};
  c2h_bits_delay_addr_REG_1 = _RAND_40[20:0];
  _RAND_41 = {1{`RANDOM}};
  REG = _RAND_41[0:0];
  _RAND_42 = {1{`RANDOM}};
  REG_1 = _RAND_42[0:0];
  _RAND_43 = {1{`RANDOM}};
  REG_2 = _RAND_43[0:0];
  _RAND_44 = {1{`RANDOM}};
  REG_3 = _RAND_44[0:0];
  _RAND_45 = {1{`RANDOM}};
  REG_4 = _RAND_45[0:0];
  _RAND_46 = {1{`RANDOM}};
  REG_5 = _RAND_46[0:0];
  _RAND_47 = {1{`RANDOM}};
  REG_6 = _RAND_47[0:0];
  _RAND_48 = {1{`RANDOM}};
  REG_7 = _RAND_48[0:0];
  _RAND_49 = {1{`RANDOM}};
  REG_8 = _RAND_49[0:0];
  _RAND_50 = {1{`RANDOM}};
  REG_9 = _RAND_50[0:0];
  _RAND_51 = {1{`RANDOM}};
  REG_10 = _RAND_51[0:0];
  _RAND_52 = {1{`RANDOM}};
  REG_11 = _RAND_52[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module RegSlice_9(
  input         clock,
  input         reset,
  output        io_upStream_ready,
  input         io_upStream_valid,
  input  [31:0] io_upStream_bits_data,
  input         io_downStream_ready,
  output        io_downStream_valid,
  output [31:0] io_downStream_bits_data
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
`endif // RANDOMIZE_REG_INIT
  reg  fwd_valid; // @[RegSlices.scala 112:34]
  reg [31:0] fwd_data_data; // @[RegSlices.scala 113:30]
  wire  fwd_ready_s = ~fwd_valid | io_downStream_ready; // @[RegSlices.scala 115:35]
  reg  bwd_ready; // @[RegSlices.scala 123:34]
  reg [31:0] bwd_data_data; // @[RegSlices.scala 124:30]
  wire  _fwd_valid_T = io_downStream_ready ? 1'h0 : fwd_valid; // @[RegSlices.scala 121:53]
  wire  bwd_valid_s = ~bwd_ready | io_upStream_valid; // @[RegSlices.scala 126:39]
  wire  _bwd_ready_T = io_upStream_valid ? 1'h0 : bwd_ready; // @[RegSlices.scala 132:53]
  assign io_upStream_ready = bwd_ready; // @[RegSlices.scala 107:31 RegSlices.scala 128:25]
  assign io_downStream_valid = fwd_valid; // @[RegSlices.scala 109:31 RegSlices.scala 116:21]
  assign io_downStream_bits_data = fwd_data_data; // @[RegSlices.scala 108:31 RegSlices.scala 117:25]
  always @(posedge clock) begin
    if (reset) begin // @[RegSlices.scala 112:34]
      fwd_valid <= 1'h0; // @[RegSlices.scala 112:34]
    end else begin
      fwd_valid <= bwd_valid_s | _fwd_valid_T; // @[RegSlices.scala 121:25]
    end
    if (fwd_ready_s) begin // @[RegSlices.scala 119:31]
      if (bwd_ready) begin // @[RegSlices.scala 127:31]
        fwd_data_data <= io_upStream_bits_data;
      end else begin
        fwd_data_data <= bwd_data_data;
      end
    end
    bwd_ready <= reset | (fwd_ready_s | _bwd_ready_T); // @[RegSlices.scala 123:34 RegSlices.scala 123:34 RegSlices.scala 132:25]
    if (bwd_ready) begin // @[RegSlices.scala 130:31]
      bwd_data_data <= io_upStream_bits_data;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  fwd_valid = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  fwd_data_data = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  bwd_ready = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  bwd_data_data = _RAND_3[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module PoorAXIL2Reg(
  input         clock,
  input         reset,
  output        io_axi_aw_ready,
  input         io_axi_aw_valid,
  input  [31:0] io_axi_aw_bits_addr,
  output        io_axi_ar_ready,
  input         io_axi_ar_valid,
  input  [31:0] io_axi_ar_bits_addr,
  output        io_axi_w_ready,
  input         io_axi_w_valid,
  input  [31:0] io_axi_w_bits_data,
  input         io_axi_r_ready,
  output        io_axi_r_valid,
  output [31:0] io_axi_r_bits_data,
  output [31:0] io_reg_control_0,
  output [31:0] io_reg_control_8,
  output [31:0] io_reg_control_9,
  output [31:0] io_reg_control_10,
  output [31:0] io_reg_control_11,
  output [31:0] io_reg_control_12,
  output [31:0] io_reg_control_13,
  output [31:0] io_reg_control_14,
  input  [31:0] io_reg_status_300,
  input  [31:0] io_reg_status_400,
  input  [31:0] io_reg_status_401,
  input  [31:0] io_reg_status_402,
  input  [31:0] io_reg_status_403,
  input  [31:0] io_reg_status_404,
  input  [31:0] io_reg_status_405,
  input  [31:0] io_reg_status_406,
  input  [31:0] io_reg_status_407,
  input  [31:0] io_reg_status_408,
  input  [31:0] io_reg_status_409,
  input  [31:0] io_reg_status_410,
  input  [31:0] io_reg_status_411,
  input  [31:0] io_reg_status_412,
  input  [31:0] io_reg_status_413,
  input  [31:0] io_reg_status_414
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
`endif // RANDOMIZE_REG_INIT
  wire  r_delay_clock; // @[PoorAXIL2Reg.scala 38:33]
  wire  r_delay_reset; // @[PoorAXIL2Reg.scala 38:33]
  wire  r_delay_io_upStream_ready; // @[PoorAXIL2Reg.scala 38:33]
  wire  r_delay_io_upStream_valid; // @[PoorAXIL2Reg.scala 38:33]
  wire [31:0] r_delay_io_upStream_bits_data; // @[PoorAXIL2Reg.scala 38:33]
  wire  r_delay_io_downStream_ready; // @[PoorAXIL2Reg.scala 38:33]
  wire  r_delay_io_downStream_valid; // @[PoorAXIL2Reg.scala 38:33]
  wire [31:0] r_delay_io_downStream_bits_data; // @[PoorAXIL2Reg.scala 38:33]
  reg [31:0] reg_control_0; // @[PoorAXIL2Reg.scala 17:30]
  reg [31:0] reg_control_8; // @[PoorAXIL2Reg.scala 17:30]
  reg [31:0] reg_control_9; // @[PoorAXIL2Reg.scala 17:30]
  reg [31:0] reg_control_10; // @[PoorAXIL2Reg.scala 17:30]
  reg [31:0] reg_control_11; // @[PoorAXIL2Reg.scala 17:30]
  reg [31:0] reg_control_12; // @[PoorAXIL2Reg.scala 17:30]
  reg [31:0] reg_control_13; // @[PoorAXIL2Reg.scala 17:30]
  reg [31:0] reg_control_14; // @[PoorAXIL2Reg.scala 17:30]
  reg [31:0] reg_status_300; // @[PoorAXIL2Reg.scala 19:29]
  reg [31:0] reg_status_400; // @[PoorAXIL2Reg.scala 19:29]
  reg [31:0] reg_status_401; // @[PoorAXIL2Reg.scala 19:29]
  reg [31:0] reg_status_402; // @[PoorAXIL2Reg.scala 19:29]
  reg [31:0] reg_status_403; // @[PoorAXIL2Reg.scala 19:29]
  reg [31:0] reg_status_404; // @[PoorAXIL2Reg.scala 19:29]
  reg [31:0] reg_status_405; // @[PoorAXIL2Reg.scala 19:29]
  reg [31:0] reg_status_406; // @[PoorAXIL2Reg.scala 19:29]
  reg [31:0] reg_status_407; // @[PoorAXIL2Reg.scala 19:29]
  reg [31:0] reg_status_408; // @[PoorAXIL2Reg.scala 19:29]
  reg [31:0] reg_status_409; // @[PoorAXIL2Reg.scala 19:29]
  reg [31:0] reg_status_410; // @[PoorAXIL2Reg.scala 19:29]
  reg [31:0] reg_status_411; // @[PoorAXIL2Reg.scala 19:29]
  reg [31:0] reg_status_412; // @[PoorAXIL2Reg.scala 19:29]
  reg [31:0] reg_status_413; // @[PoorAXIL2Reg.scala 19:29]
  reg [31:0] reg_status_414; // @[PoorAXIL2Reg.scala 19:29]
  reg  s_rd; // @[PoorAXIL2Reg.scala 30:27]
  reg  s_wr; // @[PoorAXIL2Reg.scala 31:27]
  reg [31:0] r_addr; // @[PoorAXIL2Reg.scala 41:25]
  reg [31:0] w_addr; // @[PoorAXIL2Reg.scala 42:25]
  wire  _io_axi_ar_ready_T = ~s_rd; // @[PoorAXIL2Reg.scala 44:74]
  wire [31:0] _GEN_300 = 9'h12c == r_addr[8:0] ? reg_status_300 : 32'h0; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_301 = 9'h12d == r_addr[8:0] ? 32'h0 : _GEN_300; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_302 = 9'h12e == r_addr[8:0] ? 32'h0 : _GEN_301; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_303 = 9'h12f == r_addr[8:0] ? 32'h0 : _GEN_302; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_304 = 9'h130 == r_addr[8:0] ? 32'h0 : _GEN_303; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_305 = 9'h131 == r_addr[8:0] ? 32'h0 : _GEN_304; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_306 = 9'h132 == r_addr[8:0] ? 32'h0 : _GEN_305; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_307 = 9'h133 == r_addr[8:0] ? 32'h0 : _GEN_306; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_308 = 9'h134 == r_addr[8:0] ? 32'h0 : _GEN_307; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_309 = 9'h135 == r_addr[8:0] ? 32'h0 : _GEN_308; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_310 = 9'h136 == r_addr[8:0] ? 32'h0 : _GEN_309; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_311 = 9'h137 == r_addr[8:0] ? 32'h0 : _GEN_310; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_312 = 9'h138 == r_addr[8:0] ? 32'h0 : _GEN_311; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_313 = 9'h139 == r_addr[8:0] ? 32'h0 : _GEN_312; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_314 = 9'h13a == r_addr[8:0] ? 32'h0 : _GEN_313; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_315 = 9'h13b == r_addr[8:0] ? 32'h0 : _GEN_314; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_316 = 9'h13c == r_addr[8:0] ? 32'h0 : _GEN_315; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_317 = 9'h13d == r_addr[8:0] ? 32'h0 : _GEN_316; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_318 = 9'h13e == r_addr[8:0] ? 32'h0 : _GEN_317; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_319 = 9'h13f == r_addr[8:0] ? 32'h0 : _GEN_318; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_320 = 9'h140 == r_addr[8:0] ? 32'h0 : _GEN_319; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_321 = 9'h141 == r_addr[8:0] ? 32'h0 : _GEN_320; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_322 = 9'h142 == r_addr[8:0] ? 32'h0 : _GEN_321; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_323 = 9'h143 == r_addr[8:0] ? 32'h0 : _GEN_322; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_324 = 9'h144 == r_addr[8:0] ? 32'h0 : _GEN_323; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_325 = 9'h145 == r_addr[8:0] ? 32'h0 : _GEN_324; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_326 = 9'h146 == r_addr[8:0] ? 32'h0 : _GEN_325; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_327 = 9'h147 == r_addr[8:0] ? 32'h0 : _GEN_326; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_328 = 9'h148 == r_addr[8:0] ? 32'h0 : _GEN_327; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_329 = 9'h149 == r_addr[8:0] ? 32'h0 : _GEN_328; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_330 = 9'h14a == r_addr[8:0] ? 32'h0 : _GEN_329; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_331 = 9'h14b == r_addr[8:0] ? 32'h0 : _GEN_330; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_332 = 9'h14c == r_addr[8:0] ? 32'h0 : _GEN_331; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_333 = 9'h14d == r_addr[8:0] ? 32'h0 : _GEN_332; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_334 = 9'h14e == r_addr[8:0] ? 32'h0 : _GEN_333; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_335 = 9'h14f == r_addr[8:0] ? 32'h0 : _GEN_334; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_336 = 9'h150 == r_addr[8:0] ? 32'h0 : _GEN_335; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_337 = 9'h151 == r_addr[8:0] ? 32'h0 : _GEN_336; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_338 = 9'h152 == r_addr[8:0] ? 32'h0 : _GEN_337; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_339 = 9'h153 == r_addr[8:0] ? 32'h0 : _GEN_338; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_340 = 9'h154 == r_addr[8:0] ? 32'h0 : _GEN_339; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_341 = 9'h155 == r_addr[8:0] ? 32'h0 : _GEN_340; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_342 = 9'h156 == r_addr[8:0] ? 32'h0 : _GEN_341; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_343 = 9'h157 == r_addr[8:0] ? 32'h0 : _GEN_342; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_344 = 9'h158 == r_addr[8:0] ? 32'h0 : _GEN_343; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_345 = 9'h159 == r_addr[8:0] ? 32'h0 : _GEN_344; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_346 = 9'h15a == r_addr[8:0] ? 32'h0 : _GEN_345; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_347 = 9'h15b == r_addr[8:0] ? 32'h0 : _GEN_346; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_348 = 9'h15c == r_addr[8:0] ? 32'h0 : _GEN_347; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_349 = 9'h15d == r_addr[8:0] ? 32'h0 : _GEN_348; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_350 = 9'h15e == r_addr[8:0] ? 32'h0 : _GEN_349; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_351 = 9'h15f == r_addr[8:0] ? 32'h0 : _GEN_350; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_352 = 9'h160 == r_addr[8:0] ? 32'h0 : _GEN_351; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_353 = 9'h161 == r_addr[8:0] ? 32'h0 : _GEN_352; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_354 = 9'h162 == r_addr[8:0] ? 32'h0 : _GEN_353; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_355 = 9'h163 == r_addr[8:0] ? 32'h0 : _GEN_354; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_356 = 9'h164 == r_addr[8:0] ? 32'h0 : _GEN_355; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_357 = 9'h165 == r_addr[8:0] ? 32'h0 : _GEN_356; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_358 = 9'h166 == r_addr[8:0] ? 32'h0 : _GEN_357; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_359 = 9'h167 == r_addr[8:0] ? 32'h0 : _GEN_358; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_360 = 9'h168 == r_addr[8:0] ? 32'h0 : _GEN_359; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_361 = 9'h169 == r_addr[8:0] ? 32'h0 : _GEN_360; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_362 = 9'h16a == r_addr[8:0] ? 32'h0 : _GEN_361; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_363 = 9'h16b == r_addr[8:0] ? 32'h0 : _GEN_362; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_364 = 9'h16c == r_addr[8:0] ? 32'h0 : _GEN_363; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_365 = 9'h16d == r_addr[8:0] ? 32'h0 : _GEN_364; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_366 = 9'h16e == r_addr[8:0] ? 32'h0 : _GEN_365; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_367 = 9'h16f == r_addr[8:0] ? 32'h0 : _GEN_366; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_368 = 9'h170 == r_addr[8:0] ? 32'h0 : _GEN_367; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_369 = 9'h171 == r_addr[8:0] ? 32'h0 : _GEN_368; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_370 = 9'h172 == r_addr[8:0] ? 32'h0 : _GEN_369; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_371 = 9'h173 == r_addr[8:0] ? 32'h0 : _GEN_370; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_372 = 9'h174 == r_addr[8:0] ? 32'h0 : _GEN_371; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_373 = 9'h175 == r_addr[8:0] ? 32'h0 : _GEN_372; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_374 = 9'h176 == r_addr[8:0] ? 32'h0 : _GEN_373; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_375 = 9'h177 == r_addr[8:0] ? 32'h0 : _GEN_374; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_376 = 9'h178 == r_addr[8:0] ? 32'h0 : _GEN_375; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_377 = 9'h179 == r_addr[8:0] ? 32'h0 : _GEN_376; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_378 = 9'h17a == r_addr[8:0] ? 32'h0 : _GEN_377; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_379 = 9'h17b == r_addr[8:0] ? 32'h0 : _GEN_378; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_380 = 9'h17c == r_addr[8:0] ? 32'h0 : _GEN_379; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_381 = 9'h17d == r_addr[8:0] ? 32'h0 : _GEN_380; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_382 = 9'h17e == r_addr[8:0] ? 32'h0 : _GEN_381; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_383 = 9'h17f == r_addr[8:0] ? 32'h0 : _GEN_382; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_384 = 9'h180 == r_addr[8:0] ? 32'h0 : _GEN_383; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_385 = 9'h181 == r_addr[8:0] ? 32'h0 : _GEN_384; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_386 = 9'h182 == r_addr[8:0] ? 32'h0 : _GEN_385; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_387 = 9'h183 == r_addr[8:0] ? 32'h0 : _GEN_386; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_388 = 9'h184 == r_addr[8:0] ? 32'h0 : _GEN_387; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_389 = 9'h185 == r_addr[8:0] ? 32'h0 : _GEN_388; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_390 = 9'h186 == r_addr[8:0] ? 32'h0 : _GEN_389; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_391 = 9'h187 == r_addr[8:0] ? 32'h0 : _GEN_390; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_392 = 9'h188 == r_addr[8:0] ? 32'h0 : _GEN_391; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_393 = 9'h189 == r_addr[8:0] ? 32'h0 : _GEN_392; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_394 = 9'h18a == r_addr[8:0] ? 32'h0 : _GEN_393; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_395 = 9'h18b == r_addr[8:0] ? 32'h0 : _GEN_394; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_396 = 9'h18c == r_addr[8:0] ? 32'h0 : _GEN_395; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_397 = 9'h18d == r_addr[8:0] ? 32'h0 : _GEN_396; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_398 = 9'h18e == r_addr[8:0] ? 32'h0 : _GEN_397; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_399 = 9'h18f == r_addr[8:0] ? 32'h0 : _GEN_398; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_400 = 9'h190 == r_addr[8:0] ? reg_status_400 : _GEN_399; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_401 = 9'h191 == r_addr[8:0] ? reg_status_401 : _GEN_400; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_402 = 9'h192 == r_addr[8:0] ? reg_status_402 : _GEN_401; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_403 = 9'h193 == r_addr[8:0] ? reg_status_403 : _GEN_402; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_404 = 9'h194 == r_addr[8:0] ? reg_status_404 : _GEN_403; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_405 = 9'h195 == r_addr[8:0] ? reg_status_405 : _GEN_404; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_406 = 9'h196 == r_addr[8:0] ? reg_status_406 : _GEN_405; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_407 = 9'h197 == r_addr[8:0] ? reg_status_407 : _GEN_406; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_408 = 9'h198 == r_addr[8:0] ? reg_status_408 : _GEN_407; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_409 = 9'h199 == r_addr[8:0] ? reg_status_409 : _GEN_408; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_410 = 9'h19a == r_addr[8:0] ? reg_status_410 : _GEN_409; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_411 = 9'h19b == r_addr[8:0] ? reg_status_411 : _GEN_410; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_412 = 9'h19c == r_addr[8:0] ? reg_status_412 : _GEN_411; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_413 = 9'h19d == r_addr[8:0] ? reg_status_413 : _GEN_412; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_414 = 9'h19e == r_addr[8:0] ? reg_status_414 : _GEN_413; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_415 = 9'h19f == r_addr[8:0] ? 32'h0 : _GEN_414; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_416 = 9'h1a0 == r_addr[8:0] ? 32'h0 : _GEN_415; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_417 = 9'h1a1 == r_addr[8:0] ? 32'h0 : _GEN_416; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_418 = 9'h1a2 == r_addr[8:0] ? 32'h0 : _GEN_417; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_419 = 9'h1a3 == r_addr[8:0] ? 32'h0 : _GEN_418; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_420 = 9'h1a4 == r_addr[8:0] ? 32'h0 : _GEN_419; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_421 = 9'h1a5 == r_addr[8:0] ? 32'h0 : _GEN_420; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_422 = 9'h1a6 == r_addr[8:0] ? 32'h0 : _GEN_421; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_423 = 9'h1a7 == r_addr[8:0] ? 32'h0 : _GEN_422; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_424 = 9'h1a8 == r_addr[8:0] ? 32'h0 : _GEN_423; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_425 = 9'h1a9 == r_addr[8:0] ? 32'h0 : _GEN_424; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_426 = 9'h1aa == r_addr[8:0] ? 32'h0 : _GEN_425; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_427 = 9'h1ab == r_addr[8:0] ? 32'h0 : _GEN_426; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_428 = 9'h1ac == r_addr[8:0] ? 32'h0 : _GEN_427; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_429 = 9'h1ad == r_addr[8:0] ? 32'h0 : _GEN_428; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_430 = 9'h1ae == r_addr[8:0] ? 32'h0 : _GEN_429; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_431 = 9'h1af == r_addr[8:0] ? 32'h0 : _GEN_430; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_432 = 9'h1b0 == r_addr[8:0] ? 32'h0 : _GEN_431; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_433 = 9'h1b1 == r_addr[8:0] ? 32'h0 : _GEN_432; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_434 = 9'h1b2 == r_addr[8:0] ? 32'h0 : _GEN_433; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_435 = 9'h1b3 == r_addr[8:0] ? 32'h0 : _GEN_434; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_436 = 9'h1b4 == r_addr[8:0] ? 32'h0 : _GEN_435; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_437 = 9'h1b5 == r_addr[8:0] ? 32'h0 : _GEN_436; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_438 = 9'h1b6 == r_addr[8:0] ? 32'h0 : _GEN_437; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_439 = 9'h1b7 == r_addr[8:0] ? 32'h0 : _GEN_438; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_440 = 9'h1b8 == r_addr[8:0] ? 32'h0 : _GEN_439; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_441 = 9'h1b9 == r_addr[8:0] ? 32'h0 : _GEN_440; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_442 = 9'h1ba == r_addr[8:0] ? 32'h0 : _GEN_441; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_443 = 9'h1bb == r_addr[8:0] ? 32'h0 : _GEN_442; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_444 = 9'h1bc == r_addr[8:0] ? 32'h0 : _GEN_443; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_445 = 9'h1bd == r_addr[8:0] ? 32'h0 : _GEN_444; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_446 = 9'h1be == r_addr[8:0] ? 32'h0 : _GEN_445; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_447 = 9'h1bf == r_addr[8:0] ? 32'h0 : _GEN_446; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_448 = 9'h1c0 == r_addr[8:0] ? 32'h0 : _GEN_447; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_449 = 9'h1c1 == r_addr[8:0] ? 32'h0 : _GEN_448; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_450 = 9'h1c2 == r_addr[8:0] ? 32'h0 : _GEN_449; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_451 = 9'h1c3 == r_addr[8:0] ? 32'h0 : _GEN_450; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_452 = 9'h1c4 == r_addr[8:0] ? 32'h0 : _GEN_451; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_453 = 9'h1c5 == r_addr[8:0] ? 32'h0 : _GEN_452; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_454 = 9'h1c6 == r_addr[8:0] ? 32'h0 : _GEN_453; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_455 = 9'h1c7 == r_addr[8:0] ? 32'h0 : _GEN_454; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_456 = 9'h1c8 == r_addr[8:0] ? 32'h0 : _GEN_455; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_457 = 9'h1c9 == r_addr[8:0] ? 32'h0 : _GEN_456; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_458 = 9'h1ca == r_addr[8:0] ? 32'h0 : _GEN_457; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_459 = 9'h1cb == r_addr[8:0] ? 32'h0 : _GEN_458; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_460 = 9'h1cc == r_addr[8:0] ? 32'h0 : _GEN_459; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_461 = 9'h1cd == r_addr[8:0] ? 32'h0 : _GEN_460; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_462 = 9'h1ce == r_addr[8:0] ? 32'h0 : _GEN_461; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_463 = 9'h1cf == r_addr[8:0] ? 32'h0 : _GEN_462; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_464 = 9'h1d0 == r_addr[8:0] ? 32'h0 : _GEN_463; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_465 = 9'h1d1 == r_addr[8:0] ? 32'h0 : _GEN_464; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_466 = 9'h1d2 == r_addr[8:0] ? 32'h0 : _GEN_465; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_467 = 9'h1d3 == r_addr[8:0] ? 32'h0 : _GEN_466; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_468 = 9'h1d4 == r_addr[8:0] ? 32'h0 : _GEN_467; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_469 = 9'h1d5 == r_addr[8:0] ? 32'h0 : _GEN_468; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_470 = 9'h1d6 == r_addr[8:0] ? 32'h0 : _GEN_469; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_471 = 9'h1d7 == r_addr[8:0] ? 32'h0 : _GEN_470; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_472 = 9'h1d8 == r_addr[8:0] ? 32'h0 : _GEN_471; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_473 = 9'h1d9 == r_addr[8:0] ? 32'h0 : _GEN_472; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_474 = 9'h1da == r_addr[8:0] ? 32'h0 : _GEN_473; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_475 = 9'h1db == r_addr[8:0] ? 32'h0 : _GEN_474; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_476 = 9'h1dc == r_addr[8:0] ? 32'h0 : _GEN_475; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_477 = 9'h1dd == r_addr[8:0] ? 32'h0 : _GEN_476; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_478 = 9'h1de == r_addr[8:0] ? 32'h0 : _GEN_477; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_479 = 9'h1df == r_addr[8:0] ? 32'h0 : _GEN_478; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_480 = 9'h1e0 == r_addr[8:0] ? 32'h0 : _GEN_479; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_481 = 9'h1e1 == r_addr[8:0] ? 32'h0 : _GEN_480; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_482 = 9'h1e2 == r_addr[8:0] ? 32'h0 : _GEN_481; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_483 = 9'h1e3 == r_addr[8:0] ? 32'h0 : _GEN_482; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_484 = 9'h1e4 == r_addr[8:0] ? 32'h0 : _GEN_483; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_485 = 9'h1e5 == r_addr[8:0] ? 32'h0 : _GEN_484; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_486 = 9'h1e6 == r_addr[8:0] ? 32'h0 : _GEN_485; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_487 = 9'h1e7 == r_addr[8:0] ? 32'h0 : _GEN_486; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_488 = 9'h1e8 == r_addr[8:0] ? 32'h0 : _GEN_487; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_489 = 9'h1e9 == r_addr[8:0] ? 32'h0 : _GEN_488; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_490 = 9'h1ea == r_addr[8:0] ? 32'h0 : _GEN_489; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_491 = 9'h1eb == r_addr[8:0] ? 32'h0 : _GEN_490; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_492 = 9'h1ec == r_addr[8:0] ? 32'h0 : _GEN_491; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_493 = 9'h1ed == r_addr[8:0] ? 32'h0 : _GEN_492; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_494 = 9'h1ee == r_addr[8:0] ? 32'h0 : _GEN_493; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_495 = 9'h1ef == r_addr[8:0] ? 32'h0 : _GEN_494; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_496 = 9'h1f0 == r_addr[8:0] ? 32'h0 : _GEN_495; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_497 = 9'h1f1 == r_addr[8:0] ? 32'h0 : _GEN_496; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_498 = 9'h1f2 == r_addr[8:0] ? 32'h0 : _GEN_497; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_499 = 9'h1f3 == r_addr[8:0] ? 32'h0 : _GEN_498; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_500 = 9'h1f4 == r_addr[8:0] ? 32'h0 : _GEN_499; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_501 = 9'h1f5 == r_addr[8:0] ? 32'h0 : _GEN_500; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_502 = 9'h1f6 == r_addr[8:0] ? 32'h0 : _GEN_501; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_503 = 9'h1f7 == r_addr[8:0] ? 32'h0 : _GEN_502; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_504 = 9'h1f8 == r_addr[8:0] ? 32'h0 : _GEN_503; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_505 = 9'h1f9 == r_addr[8:0] ? 32'h0 : _GEN_504; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_506 = 9'h1fa == r_addr[8:0] ? 32'h0 : _GEN_505; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_507 = 9'h1fb == r_addr[8:0] ? 32'h0 : _GEN_506; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_508 = 9'h1fc == r_addr[8:0] ? 32'h0 : _GEN_507; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_509 = 9'h1fd == r_addr[8:0] ? 32'h0 : _GEN_508; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_510 = 9'h1fe == r_addr[8:0] ? 32'h0 : _GEN_509; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire  _T_1 = io_axi_ar_ready & io_axi_ar_valid; // @[Decoupled.scala 40:37]
  wire [31:0] _r_addr_T = {{2'd0}, io_axi_ar_bits_addr[31:2]}; // @[PoorAXIL2Reg.scala 51:73]
  wire  _GEN_513 = _T_1 | s_rd; // @[PoorAXIL2Reg.scala 50:40 PoorAXIL2Reg.scala 52:57 PoorAXIL2Reg.scala 30:27]
  wire  _T_3 = r_delay_io_upStream_ready & r_delay_io_upStream_valid; // @[Decoupled.scala 40:37]
  wire  _io_axi_aw_ready_T = ~s_wr; // @[PoorAXIL2Reg.scala 62:34]
  wire  _T_4 = io_axi_w_ready & io_axi_w_valid; // @[Decoupled.scala 40:37]
  wire  _T_7 = io_axi_aw_ready & io_axi_aw_valid; // @[Decoupled.scala 40:37]
  wire [31:0] _w_addr_T = {{2'd0}, io_axi_aw_bits_addr[31:2]}; // @[PoorAXIL2Reg.scala 70:73]
  wire  _GEN_1543 = _T_7 | s_wr; // @[PoorAXIL2Reg.scala 69:40 PoorAXIL2Reg.scala 71:57 PoorAXIL2Reg.scala 31:27]
  RegSlice_9 r_delay ( // @[PoorAXIL2Reg.scala 38:33]
    .clock(r_delay_clock),
    .reset(r_delay_reset),
    .io_upStream_ready(r_delay_io_upStream_ready),
    .io_upStream_valid(r_delay_io_upStream_valid),
    .io_upStream_bits_data(r_delay_io_upStream_bits_data),
    .io_downStream_ready(r_delay_io_downStream_ready),
    .io_downStream_valid(r_delay_io_downStream_valid),
    .io_downStream_bits_data(r_delay_io_downStream_bits_data)
  );
  assign io_axi_aw_ready = ~s_wr; // @[PoorAXIL2Reg.scala 62:34]
  assign io_axi_ar_ready = ~s_rd; // @[PoorAXIL2Reg.scala 44:74]
  assign io_axi_w_ready = s_wr; // @[PoorAXIL2Reg.scala 63:34]
  assign io_axi_r_valid = r_delay_io_downStream_valid; // @[PoorAXIL2Reg.scala 47:73]
  assign io_axi_r_bits_data = r_delay_io_downStream_bits_data; // @[PoorAXIL2Reg.scala 47:73]
  assign io_reg_control_0 = reg_control_0; // @[PoorAXIL2Reg.scala 23:57]
  assign io_reg_control_8 = reg_control_8; // @[PoorAXIL2Reg.scala 23:57]
  assign io_reg_control_9 = reg_control_9; // @[PoorAXIL2Reg.scala 23:57]
  assign io_reg_control_10 = reg_control_10; // @[PoorAXIL2Reg.scala 23:57]
  assign io_reg_control_11 = reg_control_11; // @[PoorAXIL2Reg.scala 23:57]
  assign io_reg_control_12 = reg_control_12; // @[PoorAXIL2Reg.scala 23:57]
  assign io_reg_control_13 = reg_control_13; // @[PoorAXIL2Reg.scala 23:57]
  assign io_reg_control_14 = reg_control_14; // @[PoorAXIL2Reg.scala 23:57]
  assign r_delay_clock = clock;
  assign r_delay_reset = reset;
  assign r_delay_io_upStream_valid = s_rd; // @[PoorAXIL2Reg.scala 45:58]
  assign r_delay_io_upStream_bits_data = 9'h1ff == r_addr[8:0] ? 32'h0 : _GEN_510; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  assign r_delay_io_downStream_ready = io_axi_r_ready; // @[PoorAXIL2Reg.scala 47:73]
  always @(posedge clock) begin
    if (_T_4) begin // @[PoorAXIL2Reg.scala 64:23]
      if (9'h0 == w_addr[8:0]) begin // @[PoorAXIL2Reg.scala 65:41]
        reg_control_0 <= io_axi_w_bits_data; // @[PoorAXIL2Reg.scala 65:41]
      end
    end
    if (_T_4) begin // @[PoorAXIL2Reg.scala 64:23]
      if (9'h8 == w_addr[8:0]) begin // @[PoorAXIL2Reg.scala 65:41]
        reg_control_8 <= io_axi_w_bits_data; // @[PoorAXIL2Reg.scala 65:41]
      end
    end
    if (_T_4) begin // @[PoorAXIL2Reg.scala 64:23]
      if (9'h9 == w_addr[8:0]) begin // @[PoorAXIL2Reg.scala 65:41]
        reg_control_9 <= io_axi_w_bits_data; // @[PoorAXIL2Reg.scala 65:41]
      end
    end
    if (_T_4) begin // @[PoorAXIL2Reg.scala 64:23]
      if (9'ha == w_addr[8:0]) begin // @[PoorAXIL2Reg.scala 65:41]
        reg_control_10 <= io_axi_w_bits_data; // @[PoorAXIL2Reg.scala 65:41]
      end
    end
    if (_T_4) begin // @[PoorAXIL2Reg.scala 64:23]
      if (9'hb == w_addr[8:0]) begin // @[PoorAXIL2Reg.scala 65:41]
        reg_control_11 <= io_axi_w_bits_data; // @[PoorAXIL2Reg.scala 65:41]
      end
    end
    if (_T_4) begin // @[PoorAXIL2Reg.scala 64:23]
      if (9'hc == w_addr[8:0]) begin // @[PoorAXIL2Reg.scala 65:41]
        reg_control_12 <= io_axi_w_bits_data; // @[PoorAXIL2Reg.scala 65:41]
      end
    end
    if (_T_4) begin // @[PoorAXIL2Reg.scala 64:23]
      if (9'hd == w_addr[8:0]) begin // @[PoorAXIL2Reg.scala 65:41]
        reg_control_13 <= io_axi_w_bits_data; // @[PoorAXIL2Reg.scala 65:41]
      end
    end
    if (_T_4) begin // @[PoorAXIL2Reg.scala 64:23]
      if (9'he == w_addr[8:0]) begin // @[PoorAXIL2Reg.scala 65:41]
        reg_control_14 <= io_axi_w_bits_data; // @[PoorAXIL2Reg.scala 65:41]
      end
    end
    reg_status_300 <= io_reg_status_300; // @[PoorAXIL2Reg.scala 22:57]
    reg_status_400 <= io_reg_status_400; // @[PoorAXIL2Reg.scala 22:57]
    reg_status_401 <= io_reg_status_401; // @[PoorAXIL2Reg.scala 22:57]
    reg_status_402 <= io_reg_status_402; // @[PoorAXIL2Reg.scala 22:57]
    reg_status_403 <= io_reg_status_403; // @[PoorAXIL2Reg.scala 22:57]
    reg_status_404 <= io_reg_status_404; // @[PoorAXIL2Reg.scala 22:57]
    reg_status_405 <= io_reg_status_405; // @[PoorAXIL2Reg.scala 22:57]
    reg_status_406 <= io_reg_status_406; // @[PoorAXIL2Reg.scala 22:57]
    reg_status_407 <= io_reg_status_407; // @[PoorAXIL2Reg.scala 22:57]
    reg_status_408 <= io_reg_status_408; // @[PoorAXIL2Reg.scala 22:57]
    reg_status_409 <= io_reg_status_409; // @[PoorAXIL2Reg.scala 22:57]
    reg_status_410 <= io_reg_status_410; // @[PoorAXIL2Reg.scala 22:57]
    reg_status_411 <= io_reg_status_411; // @[PoorAXIL2Reg.scala 22:57]
    reg_status_412 <= io_reg_status_412; // @[PoorAXIL2Reg.scala 22:57]
    reg_status_413 <= io_reg_status_413; // @[PoorAXIL2Reg.scala 22:57]
    reg_status_414 <= io_reg_status_414; // @[PoorAXIL2Reg.scala 22:57]
    if (reset) begin // @[PoorAXIL2Reg.scala 30:27]
      s_rd <= 1'h0; // @[PoorAXIL2Reg.scala 30:27]
    end else if (_io_axi_ar_ready_T) begin // @[Conditional.scala 40:58]
      s_rd <= _GEN_513;
    end else if (s_rd) begin // @[Conditional.scala 39:67]
      if (_T_3) begin // @[PoorAXIL2Reg.scala 56:57]
        s_rd <= 1'h0; // @[PoorAXIL2Reg.scala 57:57]
      end
    end
    if (reset) begin // @[PoorAXIL2Reg.scala 31:27]
      s_wr <= 1'h0; // @[PoorAXIL2Reg.scala 31:27]
    end else if (_io_axi_aw_ready_T) begin // @[Conditional.scala 40:58]
      s_wr <= _GEN_1543;
    end else if (s_wr) begin // @[Conditional.scala 39:67]
      if (_T_4) begin // @[PoorAXIL2Reg.scala 75:39]
        s_wr <= 1'h0; // @[PoorAXIL2Reg.scala 76:57]
      end
    end
    if (_io_axi_ar_ready_T) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[PoorAXIL2Reg.scala 50:40]
        r_addr <= _r_addr_T; // @[PoorAXIL2Reg.scala 51:57]
      end
    end
    if (_io_axi_aw_ready_T) begin // @[Conditional.scala 40:58]
      if (_T_7) begin // @[PoorAXIL2Reg.scala 69:40]
        w_addr <= _w_addr_T; // @[PoorAXIL2Reg.scala 70:57]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  reg_control_0 = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  reg_control_8 = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  reg_control_9 = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  reg_control_10 = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  reg_control_11 = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  reg_control_12 = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  reg_control_13 = _RAND_6[31:0];
  _RAND_7 = {1{`RANDOM}};
  reg_control_14 = _RAND_7[31:0];
  _RAND_8 = {1{`RANDOM}};
  reg_status_300 = _RAND_8[31:0];
  _RAND_9 = {1{`RANDOM}};
  reg_status_400 = _RAND_9[31:0];
  _RAND_10 = {1{`RANDOM}};
  reg_status_401 = _RAND_10[31:0];
  _RAND_11 = {1{`RANDOM}};
  reg_status_402 = _RAND_11[31:0];
  _RAND_12 = {1{`RANDOM}};
  reg_status_403 = _RAND_12[31:0];
  _RAND_13 = {1{`RANDOM}};
  reg_status_404 = _RAND_13[31:0];
  _RAND_14 = {1{`RANDOM}};
  reg_status_405 = _RAND_14[31:0];
  _RAND_15 = {1{`RANDOM}};
  reg_status_406 = _RAND_15[31:0];
  _RAND_16 = {1{`RANDOM}};
  reg_status_407 = _RAND_16[31:0];
  _RAND_17 = {1{`RANDOM}};
  reg_status_408 = _RAND_17[31:0];
  _RAND_18 = {1{`RANDOM}};
  reg_status_409 = _RAND_18[31:0];
  _RAND_19 = {1{`RANDOM}};
  reg_status_410 = _RAND_19[31:0];
  _RAND_20 = {1{`RANDOM}};
  reg_status_411 = _RAND_20[31:0];
  _RAND_21 = {1{`RANDOM}};
  reg_status_412 = _RAND_21[31:0];
  _RAND_22 = {1{`RANDOM}};
  reg_status_413 = _RAND_22[31:0];
  _RAND_23 = {1{`RANDOM}};
  reg_status_414 = _RAND_23[31:0];
  _RAND_24 = {1{`RANDOM}};
  s_rd = _RAND_24[0:0];
  _RAND_25 = {1{`RANDOM}};
  s_wr = _RAND_25[0:0];
  _RAND_26 = {1{`RANDOM}};
  r_addr = _RAND_26[31:0];
  _RAND_27 = {1{`RANDOM}};
  w_addr = _RAND_27[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module SV_STREAM_FIFO_4(
  input          io_m_clk,
  input          io_s_clk,
  input          io_reset_n,
  input  [103:0] io_in_data,
  input          io_in_valid,
  output         io_in_ready,
  output [103:0] io_out_data,
  output         io_out_valid,
  input          io_out_ready
);
  wire [103:0] meta_m_axis_tdata; // @[Meta.scala 30:26]
  wire [12:0] meta_m_axis_tkeep; // @[Meta.scala 30:26]
  wire  meta_m_axis_tlast; // @[Meta.scala 30:26]
  wire  meta_m_axis_tvalid; // @[Meta.scala 30:26]
  wire [4:0] meta_rd_data_count_axis; // @[Meta.scala 30:26]
  wire  meta_s_axis_tready; // @[Meta.scala 30:26]
  wire [4:0] meta_wr_data_count_axis; // @[Meta.scala 30:26]
  wire  meta_m_aclk; // @[Meta.scala 30:26]
  wire  meta_m_axis_tready; // @[Meta.scala 30:26]
  wire  meta_s_aclk; // @[Meta.scala 30:26]
  wire  meta_s_aresetn; // @[Meta.scala 30:26]
  wire [103:0] meta_s_axis_tdata; // @[Meta.scala 30:26]
  wire  meta_s_axis_tdest; // @[Meta.scala 30:26]
  wire  meta_s_axis_tid; // @[Meta.scala 30:26]
  wire [12:0] meta_s_axis_tkeep; // @[Meta.scala 30:26]
  wire  meta_s_axis_tlast; // @[Meta.scala 30:26]
  wire [12:0] meta_s_axis_tstrb; // @[Meta.scala 30:26]
  wire  meta_s_axis_tuser; // @[Meta.scala 30:26]
  wire  meta_s_axis_tvalid; // @[Meta.scala 30:26]
  xpm_fifo_axis
    #(.RD_DATA_COUNT_WIDTH(5), .CLOCKING_MODE("independent_clock"), .PACKET_FIFO("false"), .USE_ADV_FEATURES("0404"), .TID_WIDTH(1), .TDEST_WIDTH(1), .PROG_EMPTY_THRESH(10), .TUSER_WIDTH(1), .FIFO_DEPTH(16), .SIM_ASSERT_CHK(0), .WR_DATA_COUNT_WIDTH(5), .ECC_MODE("no_ecc"), .FIFO_MEMORY_TYPE("auto"), .PROG_FULL_THRESH(10), .TDATA_WIDTH(104), .RELATED_CLOCKS(0), .CASCADE_HEIGHT(0), .CDC_SYNC_STAGES(2))
    meta ( // @[Meta.scala 30:26]
    .m_axis_tdata(meta_m_axis_tdata),
    .m_axis_tkeep(meta_m_axis_tkeep),
    .m_axis_tlast(meta_m_axis_tlast),
    .m_axis_tvalid(meta_m_axis_tvalid),
    .rd_data_count_axis(meta_rd_data_count_axis),
    .s_axis_tready(meta_s_axis_tready),
    .wr_data_count_axis(meta_wr_data_count_axis),
    .m_aclk(meta_m_aclk),
    .m_axis_tready(meta_m_axis_tready),
    .s_aclk(meta_s_aclk),
    .s_aresetn(meta_s_aresetn),
    .s_axis_tdata(meta_s_axis_tdata),
    .s_axis_tdest(meta_s_axis_tdest),
    .s_axis_tid(meta_s_axis_tid),
    .s_axis_tkeep(meta_s_axis_tkeep),
    .s_axis_tlast(meta_s_axis_tlast),
    .s_axis_tstrb(meta_s_axis_tstrb),
    .s_axis_tuser(meta_s_axis_tuser),
    .s_axis_tvalid(meta_s_axis_tvalid)
  );
  assign io_in_ready = meta_s_axis_tready; // @[Meta.scala 34:41]
  assign io_out_data = meta_m_axis_tdata; // @[Meta.scala 31:41]
  assign io_out_valid = meta_m_axis_tvalid; // @[Meta.scala 32:41]
  assign meta_m_aclk = io_m_clk; // @[Meta.scala 37:49]
  assign meta_m_axis_tready = io_out_ready; // @[Meta.scala 38:41]
  assign meta_s_aclk = io_s_clk; // @[Meta.scala 39:49]
  assign meta_s_aresetn = io_reset_n; // @[Meta.scala 40:49]
  assign meta_s_axis_tdata = io_in_data; // @[Meta.scala 41:41]
  assign meta_s_axis_tdest = 1'h0; // @[Meta.scala 42:41]
  assign meta_s_axis_tid = 1'h0; // @[Meta.scala 43:49]
  assign meta_s_axis_tkeep = 13'h1fff; // @[Bitwise.scala 72:12]
  assign meta_s_axis_tlast = 1'h1; // @[Meta.scala 45:41]
  assign meta_s_axis_tstrb = 13'h1fff; // @[Bitwise.scala 72:12]
  assign meta_s_axis_tuser = 1'h0; // @[Meta.scala 47:41]
  assign meta_s_axis_tvalid = io_in_valid; // @[Meta.scala 48:41]
endmodule
module XConverter_4(
  input         io_in_clk,
  input         io_out_clk,
  input         io_rstn,
  output        io_in_ready,
  input         io_in_valid,
  input  [63:0] io_in_bits_addr,
  input  [1:0]  io_in_bits_burst,
  input  [3:0]  io_in_bits_cache,
  input  [3:0]  io_in_bits_id,
  input  [7:0]  io_in_bits_len,
  input         io_in_bits_lock,
  input  [2:0]  io_in_bits_prot,
  input  [2:0]  io_in_bits_size,
  input         io_out_ready,
  output        io_out_valid,
  output [63:0] io_out_bits_addr
);
  wire  fifo_io_m_clk; // @[XConverter.scala 97:34]
  wire  fifo_io_s_clk; // @[XConverter.scala 97:34]
  wire  fifo_io_reset_n; // @[XConverter.scala 97:34]
  wire [103:0] fifo_io_in_data; // @[XConverter.scala 97:34]
  wire  fifo_io_in_valid; // @[XConverter.scala 97:34]
  wire  fifo_io_in_ready; // @[XConverter.scala 97:34]
  wire [103:0] fifo_io_out_data; // @[XConverter.scala 97:34]
  wire  fifo_io_out_valid; // @[XConverter.scala 97:34]
  wire  fifo_io_out_ready; // @[XConverter.scala 97:34]
  wire [96:0] _fifo_io_in_data_T = {io_in_bits_addr,io_in_bits_burst,io_in_bits_cache,io_in_bits_id,io_in_bits_len,
    io_in_bits_lock,io_in_bits_prot,4'h0,4'h0,io_in_bits_size}; // @[XConverter.scala 103:63]
  SV_STREAM_FIFO_4 fifo ( // @[XConverter.scala 97:34]
    .io_m_clk(fifo_io_m_clk),
    .io_s_clk(fifo_io_s_clk),
    .io_reset_n(fifo_io_reset_n),
    .io_in_data(fifo_io_in_data),
    .io_in_valid(fifo_io_in_valid),
    .io_in_ready(fifo_io_in_ready),
    .io_out_data(fifo_io_out_data),
    .io_out_valid(fifo_io_out_valid),
    .io_out_ready(fifo_io_out_ready)
  );
  assign io_in_ready = fifo_io_in_ready; // @[XConverter.scala 105:41]
  assign io_out_valid = fifo_io_out_valid; // @[XConverter.scala 108:41]
  assign io_out_bits_addr = fifo_io_out_data[96:33]; // @[XConverter.scala 107:77]
  assign fifo_io_m_clk = io_out_clk; // @[XConverter.scala 100:41]
  assign fifo_io_s_clk = io_in_clk; // @[XConverter.scala 99:41]
  assign fifo_io_reset_n = io_rstn; // @[XConverter.scala 101:41]
  assign fifo_io_in_data = {{7'd0}, _fifo_io_in_data_T}; // @[XConverter.scala 103:63]
  assign fifo_io_in_valid = io_in_valid; // @[XConverter.scala 104:41]
  assign fifo_io_out_ready = io_out_ready; // @[XConverter.scala 109:41]
endmodule
module SV_STREAM_FIFO_6(
  input          io_m_clk,
  input          io_s_clk,
  input          io_reset_n,
  input  [583:0] io_in_data,
  input          io_in_valid,
  output         io_in_ready,
  output [583:0] io_out_data,
  output         io_out_valid,
  input          io_out_ready
);
  wire [583:0] meta_m_axis_tdata; // @[Meta.scala 30:26]
  wire [72:0] meta_m_axis_tkeep; // @[Meta.scala 30:26]
  wire  meta_m_axis_tlast; // @[Meta.scala 30:26]
  wire  meta_m_axis_tvalid; // @[Meta.scala 30:26]
  wire [4:0] meta_rd_data_count_axis; // @[Meta.scala 30:26]
  wire  meta_s_axis_tready; // @[Meta.scala 30:26]
  wire [4:0] meta_wr_data_count_axis; // @[Meta.scala 30:26]
  wire  meta_m_aclk; // @[Meta.scala 30:26]
  wire  meta_m_axis_tready; // @[Meta.scala 30:26]
  wire  meta_s_aclk; // @[Meta.scala 30:26]
  wire  meta_s_aresetn; // @[Meta.scala 30:26]
  wire [583:0] meta_s_axis_tdata; // @[Meta.scala 30:26]
  wire  meta_s_axis_tdest; // @[Meta.scala 30:26]
  wire  meta_s_axis_tid; // @[Meta.scala 30:26]
  wire [72:0] meta_s_axis_tkeep; // @[Meta.scala 30:26]
  wire  meta_s_axis_tlast; // @[Meta.scala 30:26]
  wire [72:0] meta_s_axis_tstrb; // @[Meta.scala 30:26]
  wire  meta_s_axis_tuser; // @[Meta.scala 30:26]
  wire  meta_s_axis_tvalid; // @[Meta.scala 30:26]
  xpm_fifo_axis
    #(.RD_DATA_COUNT_WIDTH(5), .CLOCKING_MODE("independent_clock"), .PACKET_FIFO("false"), .USE_ADV_FEATURES("0404"), .TID_WIDTH(1), .TDEST_WIDTH(1), .PROG_EMPTY_THRESH(10), .TUSER_WIDTH(1), .FIFO_DEPTH(16), .SIM_ASSERT_CHK(0), .WR_DATA_COUNT_WIDTH(5), .ECC_MODE("no_ecc"), .FIFO_MEMORY_TYPE("auto"), .PROG_FULL_THRESH(10), .TDATA_WIDTH(584), .RELATED_CLOCKS(0), .CASCADE_HEIGHT(0), .CDC_SYNC_STAGES(2))
    meta ( // @[Meta.scala 30:26]
    .m_axis_tdata(meta_m_axis_tdata),
    .m_axis_tkeep(meta_m_axis_tkeep),
    .m_axis_tlast(meta_m_axis_tlast),
    .m_axis_tvalid(meta_m_axis_tvalid),
    .rd_data_count_axis(meta_rd_data_count_axis),
    .s_axis_tready(meta_s_axis_tready),
    .wr_data_count_axis(meta_wr_data_count_axis),
    .m_aclk(meta_m_aclk),
    .m_axis_tready(meta_m_axis_tready),
    .s_aclk(meta_s_aclk),
    .s_aresetn(meta_s_aresetn),
    .s_axis_tdata(meta_s_axis_tdata),
    .s_axis_tdest(meta_s_axis_tdest),
    .s_axis_tid(meta_s_axis_tid),
    .s_axis_tkeep(meta_s_axis_tkeep),
    .s_axis_tlast(meta_s_axis_tlast),
    .s_axis_tstrb(meta_s_axis_tstrb),
    .s_axis_tuser(meta_s_axis_tuser),
    .s_axis_tvalid(meta_s_axis_tvalid)
  );
  assign io_in_ready = meta_s_axis_tready; // @[Meta.scala 34:41]
  assign io_out_data = meta_m_axis_tdata; // @[Meta.scala 31:41]
  assign io_out_valid = meta_m_axis_tvalid; // @[Meta.scala 32:41]
  assign meta_m_aclk = io_m_clk; // @[Meta.scala 37:49]
  assign meta_m_axis_tready = io_out_ready; // @[Meta.scala 38:41]
  assign meta_s_aclk = io_s_clk; // @[Meta.scala 39:49]
  assign meta_s_aresetn = io_reset_n; // @[Meta.scala 40:49]
  assign meta_s_axis_tdata = io_in_data; // @[Meta.scala 41:41]
  assign meta_s_axis_tdest = 1'h0; // @[Meta.scala 42:41]
  assign meta_s_axis_tid = 1'h0; // @[Meta.scala 43:49]
  assign meta_s_axis_tkeep = 73'h1ffffffffffffffffff; // @[Bitwise.scala 72:12]
  assign meta_s_axis_tlast = 1'h1; // @[Meta.scala 45:41]
  assign meta_s_axis_tstrb = 73'h1ffffffffffffffffff; // @[Bitwise.scala 72:12]
  assign meta_s_axis_tuser = 1'h0; // @[Meta.scala 47:41]
  assign meta_s_axis_tvalid = io_in_valid; // @[Meta.scala 48:41]
endmodule
module XConverter_6(
  input          io_in_clk,
  input          io_out_clk,
  input          io_rstn,
  output         io_in_ready,
  input          io_in_valid,
  input  [511:0] io_in_bits_data,
  input          io_in_bits_last,
  input  [63:0]  io_in_bits_strb,
  input          io_out_ready,
  output         io_out_valid,
  output [511:0] io_out_bits_data
);
  wire  fifo_io_m_clk; // @[XConverter.scala 97:34]
  wire  fifo_io_s_clk; // @[XConverter.scala 97:34]
  wire  fifo_io_reset_n; // @[XConverter.scala 97:34]
  wire [583:0] fifo_io_in_data; // @[XConverter.scala 97:34]
  wire  fifo_io_in_valid; // @[XConverter.scala 97:34]
  wire  fifo_io_in_ready; // @[XConverter.scala 97:34]
  wire [583:0] fifo_io_out_data; // @[XConverter.scala 97:34]
  wire  fifo_io_out_valid; // @[XConverter.scala 97:34]
  wire  fifo_io_out_ready; // @[XConverter.scala 97:34]
  wire [576:0] _fifo_io_in_data_T = {io_in_bits_data,io_in_bits_last,io_in_bits_strb}; // @[XConverter.scala 103:63]
  SV_STREAM_FIFO_6 fifo ( // @[XConverter.scala 97:34]
    .io_m_clk(fifo_io_m_clk),
    .io_s_clk(fifo_io_s_clk),
    .io_reset_n(fifo_io_reset_n),
    .io_in_data(fifo_io_in_data),
    .io_in_valid(fifo_io_in_valid),
    .io_in_ready(fifo_io_in_ready),
    .io_out_data(fifo_io_out_data),
    .io_out_valid(fifo_io_out_valid),
    .io_out_ready(fifo_io_out_ready)
  );
  assign io_in_ready = fifo_io_in_ready; // @[XConverter.scala 105:41]
  assign io_out_valid = fifo_io_out_valid; // @[XConverter.scala 108:41]
  assign io_out_bits_data = fifo_io_out_data[576:65]; // @[XConverter.scala 107:77]
  assign fifo_io_m_clk = io_out_clk; // @[XConverter.scala 100:41]
  assign fifo_io_s_clk = io_in_clk; // @[XConverter.scala 99:41]
  assign fifo_io_reset_n = io_rstn; // @[XConverter.scala 101:41]
  assign fifo_io_in_data = {{7'd0}, _fifo_io_in_data_T}; // @[XConverter.scala 103:63]
  assign fifo_io_in_valid = io_in_valid; // @[XConverter.scala 104:41]
  assign fifo_io_out_ready = io_out_ready; // @[XConverter.scala 109:41]
endmodule
module SV_STREAM_FIFO_7(
  input          io_m_clk,
  input          io_s_clk,
  input          io_reset_n,
  input  [519:0] io_in_data,
  output         io_in_ready,
  output [519:0] io_out_data,
  output         io_out_valid,
  input          io_out_ready
);
  wire [519:0] meta_m_axis_tdata; // @[Meta.scala 30:26]
  wire [64:0] meta_m_axis_tkeep; // @[Meta.scala 30:26]
  wire  meta_m_axis_tlast; // @[Meta.scala 30:26]
  wire  meta_m_axis_tvalid; // @[Meta.scala 30:26]
  wire [4:0] meta_rd_data_count_axis; // @[Meta.scala 30:26]
  wire  meta_s_axis_tready; // @[Meta.scala 30:26]
  wire [4:0] meta_wr_data_count_axis; // @[Meta.scala 30:26]
  wire  meta_m_aclk; // @[Meta.scala 30:26]
  wire  meta_m_axis_tready; // @[Meta.scala 30:26]
  wire  meta_s_aclk; // @[Meta.scala 30:26]
  wire  meta_s_aresetn; // @[Meta.scala 30:26]
  wire [519:0] meta_s_axis_tdata; // @[Meta.scala 30:26]
  wire  meta_s_axis_tdest; // @[Meta.scala 30:26]
  wire  meta_s_axis_tid; // @[Meta.scala 30:26]
  wire [64:0] meta_s_axis_tkeep; // @[Meta.scala 30:26]
  wire  meta_s_axis_tlast; // @[Meta.scala 30:26]
  wire [64:0] meta_s_axis_tstrb; // @[Meta.scala 30:26]
  wire  meta_s_axis_tuser; // @[Meta.scala 30:26]
  wire  meta_s_axis_tvalid; // @[Meta.scala 30:26]
  xpm_fifo_axis
    #(.RD_DATA_COUNT_WIDTH(5), .CLOCKING_MODE("independent_clock"), .PACKET_FIFO("false"), .USE_ADV_FEATURES("0404"), .TID_WIDTH(1), .TDEST_WIDTH(1), .PROG_EMPTY_THRESH(10), .TUSER_WIDTH(1), .FIFO_DEPTH(16), .SIM_ASSERT_CHK(0), .WR_DATA_COUNT_WIDTH(5), .ECC_MODE("no_ecc"), .FIFO_MEMORY_TYPE("auto"), .PROG_FULL_THRESH(10), .TDATA_WIDTH(520), .RELATED_CLOCKS(0), .CASCADE_HEIGHT(0), .CDC_SYNC_STAGES(2))
    meta ( // @[Meta.scala 30:26]
    .m_axis_tdata(meta_m_axis_tdata),
    .m_axis_tkeep(meta_m_axis_tkeep),
    .m_axis_tlast(meta_m_axis_tlast),
    .m_axis_tvalid(meta_m_axis_tvalid),
    .rd_data_count_axis(meta_rd_data_count_axis),
    .s_axis_tready(meta_s_axis_tready),
    .wr_data_count_axis(meta_wr_data_count_axis),
    .m_aclk(meta_m_aclk),
    .m_axis_tready(meta_m_axis_tready),
    .s_aclk(meta_s_aclk),
    .s_aresetn(meta_s_aresetn),
    .s_axis_tdata(meta_s_axis_tdata),
    .s_axis_tdest(meta_s_axis_tdest),
    .s_axis_tid(meta_s_axis_tid),
    .s_axis_tkeep(meta_s_axis_tkeep),
    .s_axis_tlast(meta_s_axis_tlast),
    .s_axis_tstrb(meta_s_axis_tstrb),
    .s_axis_tuser(meta_s_axis_tuser),
    .s_axis_tvalid(meta_s_axis_tvalid)
  );
  assign io_in_ready = meta_s_axis_tready; // @[Meta.scala 34:41]
  assign io_out_data = meta_m_axis_tdata; // @[Meta.scala 31:41]
  assign io_out_valid = meta_m_axis_tvalid; // @[Meta.scala 32:41]
  assign meta_m_aclk = io_m_clk; // @[Meta.scala 37:49]
  assign meta_m_axis_tready = io_out_ready; // @[Meta.scala 38:41]
  assign meta_s_aclk = io_s_clk; // @[Meta.scala 39:49]
  assign meta_s_aresetn = io_reset_n; // @[Meta.scala 40:49]
  assign meta_s_axis_tdata = io_in_data; // @[Meta.scala 41:41]
  assign meta_s_axis_tdest = 1'h0; // @[Meta.scala 42:41]
  assign meta_s_axis_tid = 1'h0; // @[Meta.scala 43:49]
  assign meta_s_axis_tkeep = 65'h1ffffffffffffffff; // @[Bitwise.scala 72:12]
  assign meta_s_axis_tlast = 1'h1; // @[Meta.scala 45:41]
  assign meta_s_axis_tstrb = 65'h1ffffffffffffffff; // @[Bitwise.scala 72:12]
  assign meta_s_axis_tuser = 1'h0; // @[Meta.scala 47:41]
  assign meta_s_axis_tvalid = 1'h1; // @[Meta.scala 48:41]
endmodule
module XConverter_7(
  input          io_in_clk,
  input          io_out_clk,
  input          io_rstn,
  output         io_in_ready,
  input  [511:0] io_in_bits_data,
  input          io_out_ready,
  output         io_out_valid,
  output [511:0] io_out_bits_data,
  output         io_out_bits_last,
  output [1:0]   io_out_bits_resp,
  output [3:0]   io_out_bits_id
);
  wire  fifo_io_m_clk; // @[XConverter.scala 97:34]
  wire  fifo_io_s_clk; // @[XConverter.scala 97:34]
  wire  fifo_io_reset_n; // @[XConverter.scala 97:34]
  wire [519:0] fifo_io_in_data; // @[XConverter.scala 97:34]
  wire  fifo_io_in_ready; // @[XConverter.scala 97:34]
  wire [519:0] fifo_io_out_data; // @[XConverter.scala 97:34]
  wire  fifo_io_out_valid; // @[XConverter.scala 97:34]
  wire  fifo_io_out_ready; // @[XConverter.scala 97:34]
  wire [518:0] _fifo_io_in_data_T = {io_in_bits_data,1'h1,6'h0}; // @[XConverter.scala 103:63]
  SV_STREAM_FIFO_7 fifo ( // @[XConverter.scala 97:34]
    .io_m_clk(fifo_io_m_clk),
    .io_s_clk(fifo_io_s_clk),
    .io_reset_n(fifo_io_reset_n),
    .io_in_data(fifo_io_in_data),
    .io_in_ready(fifo_io_in_ready),
    .io_out_data(fifo_io_out_data),
    .io_out_valid(fifo_io_out_valid),
    .io_out_ready(fifo_io_out_ready)
  );
  assign io_in_ready = fifo_io_in_ready; // @[XConverter.scala 105:41]
  assign io_out_valid = fifo_io_out_valid; // @[XConverter.scala 108:41]
  assign io_out_bits_data = fifo_io_out_data[518:7]; // @[XConverter.scala 107:77]
  assign io_out_bits_last = fifo_io_out_data[6]; // @[XConverter.scala 107:77]
  assign io_out_bits_resp = fifo_io_out_data[5:4]; // @[XConverter.scala 107:77]
  assign io_out_bits_id = fifo_io_out_data[3:0]; // @[XConverter.scala 107:77]
  assign fifo_io_m_clk = io_out_clk; // @[XConverter.scala 100:41]
  assign fifo_io_s_clk = io_in_clk; // @[XConverter.scala 99:41]
  assign fifo_io_reset_n = io_rstn; // @[XConverter.scala 101:41]
  assign fifo_io_in_data = {{1'd0}, _fifo_io_in_data_T}; // @[XConverter.scala 103:63]
  assign fifo_io_out_ready = io_out_ready; // @[XConverter.scala 109:41]
endmodule
module SV_STREAM_FIFO_8(
  input        io_m_clk,
  input        io_s_clk,
  input        io_reset_n,
  output [7:0] io_out_data,
  output       io_out_valid,
  input        io_out_ready
);
  wire [7:0] meta_m_axis_tdata; // @[Meta.scala 30:26]
  wire  meta_m_axis_tkeep; // @[Meta.scala 30:26]
  wire  meta_m_axis_tlast; // @[Meta.scala 30:26]
  wire  meta_m_axis_tvalid; // @[Meta.scala 30:26]
  wire [4:0] meta_rd_data_count_axis; // @[Meta.scala 30:26]
  wire  meta_s_axis_tready; // @[Meta.scala 30:26]
  wire [4:0] meta_wr_data_count_axis; // @[Meta.scala 30:26]
  wire  meta_m_aclk; // @[Meta.scala 30:26]
  wire  meta_m_axis_tready; // @[Meta.scala 30:26]
  wire  meta_s_aclk; // @[Meta.scala 30:26]
  wire  meta_s_aresetn; // @[Meta.scala 30:26]
  wire [7:0] meta_s_axis_tdata; // @[Meta.scala 30:26]
  wire  meta_s_axis_tdest; // @[Meta.scala 30:26]
  wire  meta_s_axis_tid; // @[Meta.scala 30:26]
  wire  meta_s_axis_tkeep; // @[Meta.scala 30:26]
  wire  meta_s_axis_tlast; // @[Meta.scala 30:26]
  wire  meta_s_axis_tstrb; // @[Meta.scala 30:26]
  wire  meta_s_axis_tuser; // @[Meta.scala 30:26]
  wire  meta_s_axis_tvalid; // @[Meta.scala 30:26]
  xpm_fifo_axis
    #(.RD_DATA_COUNT_WIDTH(5), .CLOCKING_MODE("independent_clock"), .PACKET_FIFO("false"), .USE_ADV_FEATURES("0404"), .TID_WIDTH(1), .TDEST_WIDTH(1), .PROG_EMPTY_THRESH(10), .TUSER_WIDTH(1), .FIFO_DEPTH(16), .SIM_ASSERT_CHK(0), .WR_DATA_COUNT_WIDTH(5), .ECC_MODE("no_ecc"), .FIFO_MEMORY_TYPE("auto"), .PROG_FULL_THRESH(10), .TDATA_WIDTH(8), .RELATED_CLOCKS(0), .CASCADE_HEIGHT(0), .CDC_SYNC_STAGES(2))
    meta ( // @[Meta.scala 30:26]
    .m_axis_tdata(meta_m_axis_tdata),
    .m_axis_tkeep(meta_m_axis_tkeep),
    .m_axis_tlast(meta_m_axis_tlast),
    .m_axis_tvalid(meta_m_axis_tvalid),
    .rd_data_count_axis(meta_rd_data_count_axis),
    .s_axis_tready(meta_s_axis_tready),
    .wr_data_count_axis(meta_wr_data_count_axis),
    .m_aclk(meta_m_aclk),
    .m_axis_tready(meta_m_axis_tready),
    .s_aclk(meta_s_aclk),
    .s_aresetn(meta_s_aresetn),
    .s_axis_tdata(meta_s_axis_tdata),
    .s_axis_tdest(meta_s_axis_tdest),
    .s_axis_tid(meta_s_axis_tid),
    .s_axis_tkeep(meta_s_axis_tkeep),
    .s_axis_tlast(meta_s_axis_tlast),
    .s_axis_tstrb(meta_s_axis_tstrb),
    .s_axis_tuser(meta_s_axis_tuser),
    .s_axis_tvalid(meta_s_axis_tvalid)
  );
  assign io_out_data = meta_m_axis_tdata; // @[Meta.scala 31:41]
  assign io_out_valid = meta_m_axis_tvalid; // @[Meta.scala 32:41]
  assign meta_m_aclk = io_m_clk; // @[Meta.scala 37:49]
  assign meta_m_axis_tready = io_out_ready; // @[Meta.scala 38:41]
  assign meta_s_aclk = io_s_clk; // @[Meta.scala 39:49]
  assign meta_s_aresetn = io_reset_n; // @[Meta.scala 40:49]
  assign meta_s_axis_tdata = 8'h0; // @[Meta.scala 41:41]
  assign meta_s_axis_tdest = 1'h0; // @[Meta.scala 42:41]
  assign meta_s_axis_tid = 1'h0; // @[Meta.scala 43:49]
  assign meta_s_axis_tkeep = 1'h1; // @[Meta.scala 44:41]
  assign meta_s_axis_tlast = 1'h1; // @[Meta.scala 45:41]
  assign meta_s_axis_tstrb = 1'h1; // @[Meta.scala 46:41]
  assign meta_s_axis_tuser = 1'h0; // @[Meta.scala 47:41]
  assign meta_s_axis_tvalid = 1'h1; // @[Meta.scala 48:41]
endmodule
module XConverter_8(
  input        io_in_clk,
  input        io_out_clk,
  input        io_rstn,
  input        io_out_ready,
  output       io_out_valid,
  output [3:0] io_out_bits_id,
  output [1:0] io_out_bits_resp
);
  wire  fifo_io_m_clk; // @[XConverter.scala 97:34]
  wire  fifo_io_s_clk; // @[XConverter.scala 97:34]
  wire  fifo_io_reset_n; // @[XConverter.scala 97:34]
  wire [7:0] fifo_io_out_data; // @[XConverter.scala 97:34]
  wire  fifo_io_out_valid; // @[XConverter.scala 97:34]
  wire  fifo_io_out_ready; // @[XConverter.scala 97:34]
  SV_STREAM_FIFO_8 fifo ( // @[XConverter.scala 97:34]
    .io_m_clk(fifo_io_m_clk),
    .io_s_clk(fifo_io_s_clk),
    .io_reset_n(fifo_io_reset_n),
    .io_out_data(fifo_io_out_data),
    .io_out_valid(fifo_io_out_valid),
    .io_out_ready(fifo_io_out_ready)
  );
  assign io_out_valid = fifo_io_out_valid; // @[XConverter.scala 108:41]
  assign io_out_bits_id = fifo_io_out_data[5:2]; // @[XConverter.scala 107:77]
  assign io_out_bits_resp = fifo_io_out_data[1:0]; // @[XConverter.scala 107:77]
  assign fifo_io_m_clk = io_out_clk; // @[XConverter.scala 100:41]
  assign fifo_io_s_clk = io_in_clk; // @[XConverter.scala 99:41]
  assign fifo_io_reset_n = io_rstn; // @[XConverter.scala 101:41]
  assign fifo_io_out_ready = io_out_ready; // @[XConverter.scala 109:41]
endmodule
module SV_STREAM_FIFO_9(
  input         io_m_clk,
  input         io_s_clk,
  input         io_reset_n,
  input  [55:0] io_in_data,
  input         io_in_valid,
  output        io_in_ready,
  output [55:0] io_out_data,
  output        io_out_valid,
  input         io_out_ready
);
  wire [55:0] meta_m_axis_tdata; // @[Meta.scala 30:26]
  wire [6:0] meta_m_axis_tkeep; // @[Meta.scala 30:26]
  wire  meta_m_axis_tlast; // @[Meta.scala 30:26]
  wire  meta_m_axis_tvalid; // @[Meta.scala 30:26]
  wire [4:0] meta_rd_data_count_axis; // @[Meta.scala 30:26]
  wire  meta_s_axis_tready; // @[Meta.scala 30:26]
  wire [4:0] meta_wr_data_count_axis; // @[Meta.scala 30:26]
  wire  meta_m_aclk; // @[Meta.scala 30:26]
  wire  meta_m_axis_tready; // @[Meta.scala 30:26]
  wire  meta_s_aclk; // @[Meta.scala 30:26]
  wire  meta_s_aresetn; // @[Meta.scala 30:26]
  wire [55:0] meta_s_axis_tdata; // @[Meta.scala 30:26]
  wire  meta_s_axis_tdest; // @[Meta.scala 30:26]
  wire  meta_s_axis_tid; // @[Meta.scala 30:26]
  wire [6:0] meta_s_axis_tkeep; // @[Meta.scala 30:26]
  wire  meta_s_axis_tlast; // @[Meta.scala 30:26]
  wire [6:0] meta_s_axis_tstrb; // @[Meta.scala 30:26]
  wire  meta_s_axis_tuser; // @[Meta.scala 30:26]
  wire  meta_s_axis_tvalid; // @[Meta.scala 30:26]
  xpm_fifo_axis
    #(.RD_DATA_COUNT_WIDTH(5), .CLOCKING_MODE("independent_clock"), .PACKET_FIFO("false"), .USE_ADV_FEATURES("0404"), .TID_WIDTH(1), .TDEST_WIDTH(1), .PROG_EMPTY_THRESH(10), .TUSER_WIDTH(1), .FIFO_DEPTH(16), .SIM_ASSERT_CHK(0), .WR_DATA_COUNT_WIDTH(5), .ECC_MODE("no_ecc"), .FIFO_MEMORY_TYPE("auto"), .PROG_FULL_THRESH(10), .TDATA_WIDTH(56), .RELATED_CLOCKS(0), .CASCADE_HEIGHT(0), .CDC_SYNC_STAGES(2))
    meta ( // @[Meta.scala 30:26]
    .m_axis_tdata(meta_m_axis_tdata),
    .m_axis_tkeep(meta_m_axis_tkeep),
    .m_axis_tlast(meta_m_axis_tlast),
    .m_axis_tvalid(meta_m_axis_tvalid),
    .rd_data_count_axis(meta_rd_data_count_axis),
    .s_axis_tready(meta_s_axis_tready),
    .wr_data_count_axis(meta_wr_data_count_axis),
    .m_aclk(meta_m_aclk),
    .m_axis_tready(meta_m_axis_tready),
    .s_aclk(meta_s_aclk),
    .s_aresetn(meta_s_aresetn),
    .s_axis_tdata(meta_s_axis_tdata),
    .s_axis_tdest(meta_s_axis_tdest),
    .s_axis_tid(meta_s_axis_tid),
    .s_axis_tkeep(meta_s_axis_tkeep),
    .s_axis_tlast(meta_s_axis_tlast),
    .s_axis_tstrb(meta_s_axis_tstrb),
    .s_axis_tuser(meta_s_axis_tuser),
    .s_axis_tvalid(meta_s_axis_tvalid)
  );
  assign io_in_ready = meta_s_axis_tready; // @[Meta.scala 34:41]
  assign io_out_data = meta_m_axis_tdata; // @[Meta.scala 31:41]
  assign io_out_valid = meta_m_axis_tvalid; // @[Meta.scala 32:41]
  assign meta_m_aclk = io_m_clk; // @[Meta.scala 37:49]
  assign meta_m_axis_tready = io_out_ready; // @[Meta.scala 38:41]
  assign meta_s_aclk = io_s_clk; // @[Meta.scala 39:49]
  assign meta_s_aresetn = io_reset_n; // @[Meta.scala 40:49]
  assign meta_s_axis_tdata = io_in_data; // @[Meta.scala 41:41]
  assign meta_s_axis_tdest = 1'h0; // @[Meta.scala 42:41]
  assign meta_s_axis_tid = 1'h0; // @[Meta.scala 43:49]
  assign meta_s_axis_tkeep = 7'h7f; // @[Bitwise.scala 72:12]
  assign meta_s_axis_tlast = 1'h1; // @[Meta.scala 45:41]
  assign meta_s_axis_tstrb = 7'h7f; // @[Bitwise.scala 72:12]
  assign meta_s_axis_tuser = 1'h0; // @[Meta.scala 47:41]
  assign meta_s_axis_tvalid = io_in_valid; // @[Meta.scala 48:41]
endmodule
module XConverter_9(
  input         io_in_clk,
  input         io_out_clk,
  input         io_rstn,
  output        io_in_ready,
  input         io_in_valid,
  input  [31:0] io_in_bits_addr,
  input         io_out_ready,
  output        io_out_valid,
  output [31:0] io_out_bits_addr
);
  wire  fifo_io_m_clk; // @[XConverter.scala 97:34]
  wire  fifo_io_s_clk; // @[XConverter.scala 97:34]
  wire  fifo_io_reset_n; // @[XConverter.scala 97:34]
  wire [55:0] fifo_io_in_data; // @[XConverter.scala 97:34]
  wire  fifo_io_in_valid; // @[XConverter.scala 97:34]
  wire  fifo_io_in_ready; // @[XConverter.scala 97:34]
  wire [55:0] fifo_io_out_data; // @[XConverter.scala 97:34]
  wire  fifo_io_out_valid; // @[XConverter.scala 97:34]
  wire  fifo_io_out_ready; // @[XConverter.scala 97:34]
  wire [52:0] _fifo_io_in_data_T = {io_in_bits_addr,2'h0,4'h0,1'h0,14'h0}; // @[XConverter.scala 103:63]
  SV_STREAM_FIFO_9 fifo ( // @[XConverter.scala 97:34]
    .io_m_clk(fifo_io_m_clk),
    .io_s_clk(fifo_io_s_clk),
    .io_reset_n(fifo_io_reset_n),
    .io_in_data(fifo_io_in_data),
    .io_in_valid(fifo_io_in_valid),
    .io_in_ready(fifo_io_in_ready),
    .io_out_data(fifo_io_out_data),
    .io_out_valid(fifo_io_out_valid),
    .io_out_ready(fifo_io_out_ready)
  );
  assign io_in_ready = fifo_io_in_ready; // @[XConverter.scala 105:41]
  assign io_out_valid = fifo_io_out_valid; // @[XConverter.scala 108:41]
  assign io_out_bits_addr = fifo_io_out_data[52:21]; // @[XConverter.scala 107:77]
  assign fifo_io_m_clk = io_out_clk; // @[XConverter.scala 100:41]
  assign fifo_io_s_clk = io_in_clk; // @[XConverter.scala 99:41]
  assign fifo_io_reset_n = io_rstn; // @[XConverter.scala 101:41]
  assign fifo_io_in_data = {{3'd0}, _fifo_io_in_data_T}; // @[XConverter.scala 103:63]
  assign fifo_io_in_valid = io_in_valid; // @[XConverter.scala 104:41]
  assign fifo_io_out_ready = io_out_ready; // @[XConverter.scala 109:41]
endmodule
module SV_STREAM_FIFO_11(
  input         io_m_clk,
  input         io_s_clk,
  input         io_reset_n,
  input  [39:0] io_in_data,
  input         io_in_valid,
  output        io_in_ready,
  output [39:0] io_out_data,
  output        io_out_valid,
  input         io_out_ready
);
  wire [39:0] meta_m_axis_tdata; // @[Meta.scala 30:26]
  wire [4:0] meta_m_axis_tkeep; // @[Meta.scala 30:26]
  wire  meta_m_axis_tlast; // @[Meta.scala 30:26]
  wire  meta_m_axis_tvalid; // @[Meta.scala 30:26]
  wire [4:0] meta_rd_data_count_axis; // @[Meta.scala 30:26]
  wire  meta_s_axis_tready; // @[Meta.scala 30:26]
  wire [4:0] meta_wr_data_count_axis; // @[Meta.scala 30:26]
  wire  meta_m_aclk; // @[Meta.scala 30:26]
  wire  meta_m_axis_tready; // @[Meta.scala 30:26]
  wire  meta_s_aclk; // @[Meta.scala 30:26]
  wire  meta_s_aresetn; // @[Meta.scala 30:26]
  wire [39:0] meta_s_axis_tdata; // @[Meta.scala 30:26]
  wire  meta_s_axis_tdest; // @[Meta.scala 30:26]
  wire  meta_s_axis_tid; // @[Meta.scala 30:26]
  wire [4:0] meta_s_axis_tkeep; // @[Meta.scala 30:26]
  wire  meta_s_axis_tlast; // @[Meta.scala 30:26]
  wire [4:0] meta_s_axis_tstrb; // @[Meta.scala 30:26]
  wire  meta_s_axis_tuser; // @[Meta.scala 30:26]
  wire  meta_s_axis_tvalid; // @[Meta.scala 30:26]
  xpm_fifo_axis
    #(.RD_DATA_COUNT_WIDTH(5), .CLOCKING_MODE("independent_clock"), .PACKET_FIFO("false"), .USE_ADV_FEATURES("0404"), .TID_WIDTH(1), .TDEST_WIDTH(1), .PROG_EMPTY_THRESH(10), .TUSER_WIDTH(1), .FIFO_DEPTH(16), .SIM_ASSERT_CHK(0), .WR_DATA_COUNT_WIDTH(5), .ECC_MODE("no_ecc"), .FIFO_MEMORY_TYPE("auto"), .PROG_FULL_THRESH(10), .TDATA_WIDTH(40), .RELATED_CLOCKS(0), .CASCADE_HEIGHT(0), .CDC_SYNC_STAGES(2))
    meta ( // @[Meta.scala 30:26]
    .m_axis_tdata(meta_m_axis_tdata),
    .m_axis_tkeep(meta_m_axis_tkeep),
    .m_axis_tlast(meta_m_axis_tlast),
    .m_axis_tvalid(meta_m_axis_tvalid),
    .rd_data_count_axis(meta_rd_data_count_axis),
    .s_axis_tready(meta_s_axis_tready),
    .wr_data_count_axis(meta_wr_data_count_axis),
    .m_aclk(meta_m_aclk),
    .m_axis_tready(meta_m_axis_tready),
    .s_aclk(meta_s_aclk),
    .s_aresetn(meta_s_aresetn),
    .s_axis_tdata(meta_s_axis_tdata),
    .s_axis_tdest(meta_s_axis_tdest),
    .s_axis_tid(meta_s_axis_tid),
    .s_axis_tkeep(meta_s_axis_tkeep),
    .s_axis_tlast(meta_s_axis_tlast),
    .s_axis_tstrb(meta_s_axis_tstrb),
    .s_axis_tuser(meta_s_axis_tuser),
    .s_axis_tvalid(meta_s_axis_tvalid)
  );
  assign io_in_ready = meta_s_axis_tready; // @[Meta.scala 34:41]
  assign io_out_data = meta_m_axis_tdata; // @[Meta.scala 31:41]
  assign io_out_valid = meta_m_axis_tvalid; // @[Meta.scala 32:41]
  assign meta_m_aclk = io_m_clk; // @[Meta.scala 37:49]
  assign meta_m_axis_tready = io_out_ready; // @[Meta.scala 38:41]
  assign meta_s_aclk = io_s_clk; // @[Meta.scala 39:49]
  assign meta_s_aresetn = io_reset_n; // @[Meta.scala 40:49]
  assign meta_s_axis_tdata = io_in_data; // @[Meta.scala 41:41]
  assign meta_s_axis_tdest = 1'h0; // @[Meta.scala 42:41]
  assign meta_s_axis_tid = 1'h0; // @[Meta.scala 43:49]
  assign meta_s_axis_tkeep = 5'h1f; // @[Bitwise.scala 72:12]
  assign meta_s_axis_tlast = 1'h1; // @[Meta.scala 45:41]
  assign meta_s_axis_tstrb = 5'h1f; // @[Bitwise.scala 72:12]
  assign meta_s_axis_tuser = 1'h0; // @[Meta.scala 47:41]
  assign meta_s_axis_tvalid = io_in_valid; // @[Meta.scala 48:41]
endmodule
module XConverter_11(
  input         io_in_clk,
  input         io_out_clk,
  input         io_rstn,
  output        io_in_ready,
  input         io_in_valid,
  input  [31:0] io_in_bits_data,
  input  [3:0]  io_in_bits_strb,
  input         io_out_ready,
  output        io_out_valid,
  output [31:0] io_out_bits_data
);
  wire  fifo_io_m_clk; // @[XConverter.scala 97:34]
  wire  fifo_io_s_clk; // @[XConverter.scala 97:34]
  wire  fifo_io_reset_n; // @[XConverter.scala 97:34]
  wire [39:0] fifo_io_in_data; // @[XConverter.scala 97:34]
  wire  fifo_io_in_valid; // @[XConverter.scala 97:34]
  wire  fifo_io_in_ready; // @[XConverter.scala 97:34]
  wire [39:0] fifo_io_out_data; // @[XConverter.scala 97:34]
  wire  fifo_io_out_valid; // @[XConverter.scala 97:34]
  wire  fifo_io_out_ready; // @[XConverter.scala 97:34]
  wire [36:0] _fifo_io_in_data_T = {io_in_bits_data,1'h1,io_in_bits_strb}; // @[XConverter.scala 103:63]
  SV_STREAM_FIFO_11 fifo ( // @[XConverter.scala 97:34]
    .io_m_clk(fifo_io_m_clk),
    .io_s_clk(fifo_io_s_clk),
    .io_reset_n(fifo_io_reset_n),
    .io_in_data(fifo_io_in_data),
    .io_in_valid(fifo_io_in_valid),
    .io_in_ready(fifo_io_in_ready),
    .io_out_data(fifo_io_out_data),
    .io_out_valid(fifo_io_out_valid),
    .io_out_ready(fifo_io_out_ready)
  );
  assign io_in_ready = fifo_io_in_ready; // @[XConverter.scala 105:41]
  assign io_out_valid = fifo_io_out_valid; // @[XConverter.scala 108:41]
  assign io_out_bits_data = fifo_io_out_data[36:5]; // @[XConverter.scala 107:77]
  assign fifo_io_m_clk = io_out_clk; // @[XConverter.scala 100:41]
  assign fifo_io_s_clk = io_in_clk; // @[XConverter.scala 99:41]
  assign fifo_io_reset_n = io_rstn; // @[XConverter.scala 101:41]
  assign fifo_io_in_data = {{3'd0}, _fifo_io_in_data_T}; // @[XConverter.scala 103:63]
  assign fifo_io_in_valid = io_in_valid; // @[XConverter.scala 104:41]
  assign fifo_io_out_ready = io_out_ready; // @[XConverter.scala 109:41]
endmodule
module XConverter_12(
  input         io_in_clk,
  input         io_out_clk,
  input         io_rstn,
  output        io_in_ready,
  input         io_in_valid,
  input  [31:0] io_in_bits_data,
  input         io_out_ready,
  output        io_out_valid,
  output [31:0] io_out_bits_data,
  output [1:0]  io_out_bits_resp
);
  wire  fifo_io_m_clk; // @[XConverter.scala 97:34]
  wire  fifo_io_s_clk; // @[XConverter.scala 97:34]
  wire  fifo_io_reset_n; // @[XConverter.scala 97:34]
  wire [39:0] fifo_io_in_data; // @[XConverter.scala 97:34]
  wire  fifo_io_in_valid; // @[XConverter.scala 97:34]
  wire  fifo_io_in_ready; // @[XConverter.scala 97:34]
  wire [39:0] fifo_io_out_data; // @[XConverter.scala 97:34]
  wire  fifo_io_out_valid; // @[XConverter.scala 97:34]
  wire  fifo_io_out_ready; // @[XConverter.scala 97:34]
  wire [34:0] _fifo_io_in_data_T = {io_in_bits_data,1'h0,2'h0}; // @[XConverter.scala 103:63]
  SV_STREAM_FIFO_11 fifo ( // @[XConverter.scala 97:34]
    .io_m_clk(fifo_io_m_clk),
    .io_s_clk(fifo_io_s_clk),
    .io_reset_n(fifo_io_reset_n),
    .io_in_data(fifo_io_in_data),
    .io_in_valid(fifo_io_in_valid),
    .io_in_ready(fifo_io_in_ready),
    .io_out_data(fifo_io_out_data),
    .io_out_valid(fifo_io_out_valid),
    .io_out_ready(fifo_io_out_ready)
  );
  assign io_in_ready = fifo_io_in_ready; // @[XConverter.scala 105:41]
  assign io_out_valid = fifo_io_out_valid; // @[XConverter.scala 108:41]
  assign io_out_bits_data = fifo_io_out_data[34:3]; // @[XConverter.scala 107:77]
  assign io_out_bits_resp = fifo_io_out_data[1:0]; // @[XConverter.scala 107:77]
  assign fifo_io_m_clk = io_out_clk; // @[XConverter.scala 100:41]
  assign fifo_io_s_clk = io_in_clk; // @[XConverter.scala 99:41]
  assign fifo_io_reset_n = io_rstn; // @[XConverter.scala 101:41]
  assign fifo_io_in_data = {{5'd0}, _fifo_io_in_data_T}; // @[XConverter.scala 103:63]
  assign fifo_io_in_valid = io_in_valid; // @[XConverter.scala 104:41]
  assign fifo_io_out_ready = io_out_ready; // @[XConverter.scala 109:41]
endmodule
module XConverter_13(
  input        io_in_clk,
  input        io_out_clk,
  input        io_rstn,
  input        io_out_ready,
  output       io_out_valid,
  output [1:0] io_out_bits_resp
);
  wire  fifo_io_m_clk; // @[XConverter.scala 97:34]
  wire  fifo_io_s_clk; // @[XConverter.scala 97:34]
  wire  fifo_io_reset_n; // @[XConverter.scala 97:34]
  wire [7:0] fifo_io_out_data; // @[XConverter.scala 97:34]
  wire  fifo_io_out_valid; // @[XConverter.scala 97:34]
  wire  fifo_io_out_ready; // @[XConverter.scala 97:34]
  SV_STREAM_FIFO_8 fifo ( // @[XConverter.scala 97:34]
    .io_m_clk(fifo_io_m_clk),
    .io_s_clk(fifo_io_s_clk),
    .io_reset_n(fifo_io_reset_n),
    .io_out_data(fifo_io_out_data),
    .io_out_valid(fifo_io_out_valid),
    .io_out_ready(fifo_io_out_ready)
  );
  assign io_out_valid = fifo_io_out_valid; // @[XConverter.scala 108:41]
  assign io_out_bits_resp = fifo_io_out_data[1:0]; // @[XConverter.scala 107:77]
  assign fifo_io_m_clk = io_out_clk; // @[XConverter.scala 100:41]
  assign fifo_io_s_clk = io_in_clk; // @[XConverter.scala 99:41]
  assign fifo_io_reset_n = io_rstn; // @[XConverter.scala 101:41]
  assign fifo_io_out_ready = io_out_ready; // @[XConverter.scala 109:41]
endmodule
module Queue_2(
  input          clock,
  input          reset,
  input          io_deq_ready,
  output         io_deq_valid,
  output [511:0] io_deq_bits_data,
  output [31:0]  io_deq_bits_tcrc,
  output         io_deq_bits_ctrl_marker,
  output [6:0]   io_deq_bits_ctrl_ecc,
  output [31:0]  io_deq_bits_ctrl_len,
  output [2:0]   io_deq_bits_ctrl_port_id,
  output [10:0]  io_deq_bits_ctrl_qid,
  output         io_deq_bits_ctrl_has_cmpt,
  output         io_deq_bits_last,
  output [5:0]   io_deq_bits_mty
);
`ifdef RANDOMIZE_MEM_INIT
  reg [511:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_10;
`endif // RANDOMIZE_REG_INIT
  reg [511:0] ram_data [0:15]; // @[Decoupled.scala 218:16]
  wire [511:0] ram_data_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16]
  wire [3:0] ram_data_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16]
  wire [511:0] ram_data_MPORT_data; // @[Decoupled.scala 218:16]
  wire [3:0] ram_data_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_data_MPORT_mask; // @[Decoupled.scala 218:16]
  wire  ram_data_MPORT_en; // @[Decoupled.scala 218:16]
  reg [31:0] ram_tcrc [0:15]; // @[Decoupled.scala 218:16]
  wire [31:0] ram_tcrc_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16]
  wire [3:0] ram_tcrc_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16]
  wire [31:0] ram_tcrc_MPORT_data; // @[Decoupled.scala 218:16]
  wire [3:0] ram_tcrc_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_tcrc_MPORT_mask; // @[Decoupled.scala 218:16]
  wire  ram_tcrc_MPORT_en; // @[Decoupled.scala 218:16]
  reg  ram_ctrl_marker [0:15]; // @[Decoupled.scala 218:16]
  wire  ram_ctrl_marker_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16]
  wire [3:0] ram_ctrl_marker_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_ctrl_marker_MPORT_data; // @[Decoupled.scala 218:16]
  wire [3:0] ram_ctrl_marker_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_ctrl_marker_MPORT_mask; // @[Decoupled.scala 218:16]
  wire  ram_ctrl_marker_MPORT_en; // @[Decoupled.scala 218:16]
  reg [6:0] ram_ctrl_ecc [0:15]; // @[Decoupled.scala 218:16]
  wire [6:0] ram_ctrl_ecc_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16]
  wire [3:0] ram_ctrl_ecc_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16]
  wire [6:0] ram_ctrl_ecc_MPORT_data; // @[Decoupled.scala 218:16]
  wire [3:0] ram_ctrl_ecc_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_ctrl_ecc_MPORT_mask; // @[Decoupled.scala 218:16]
  wire  ram_ctrl_ecc_MPORT_en; // @[Decoupled.scala 218:16]
  reg [31:0] ram_ctrl_len [0:15]; // @[Decoupled.scala 218:16]
  wire [31:0] ram_ctrl_len_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16]
  wire [3:0] ram_ctrl_len_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16]
  wire [31:0] ram_ctrl_len_MPORT_data; // @[Decoupled.scala 218:16]
  wire [3:0] ram_ctrl_len_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_ctrl_len_MPORT_mask; // @[Decoupled.scala 218:16]
  wire  ram_ctrl_len_MPORT_en; // @[Decoupled.scala 218:16]
  reg [2:0] ram_ctrl_port_id [0:15]; // @[Decoupled.scala 218:16]
  wire [2:0] ram_ctrl_port_id_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16]
  wire [3:0] ram_ctrl_port_id_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16]
  wire [2:0] ram_ctrl_port_id_MPORT_data; // @[Decoupled.scala 218:16]
  wire [3:0] ram_ctrl_port_id_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_ctrl_port_id_MPORT_mask; // @[Decoupled.scala 218:16]
  wire  ram_ctrl_port_id_MPORT_en; // @[Decoupled.scala 218:16]
  reg [10:0] ram_ctrl_qid [0:15]; // @[Decoupled.scala 218:16]
  wire [10:0] ram_ctrl_qid_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16]
  wire [3:0] ram_ctrl_qid_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16]
  wire [10:0] ram_ctrl_qid_MPORT_data; // @[Decoupled.scala 218:16]
  wire [3:0] ram_ctrl_qid_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_ctrl_qid_MPORT_mask; // @[Decoupled.scala 218:16]
  wire  ram_ctrl_qid_MPORT_en; // @[Decoupled.scala 218:16]
  reg  ram_ctrl_has_cmpt [0:15]; // @[Decoupled.scala 218:16]
  wire  ram_ctrl_has_cmpt_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16]
  wire [3:0] ram_ctrl_has_cmpt_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_ctrl_has_cmpt_MPORT_data; // @[Decoupled.scala 218:16]
  wire [3:0] ram_ctrl_has_cmpt_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_ctrl_has_cmpt_MPORT_mask; // @[Decoupled.scala 218:16]
  wire  ram_ctrl_has_cmpt_MPORT_en; // @[Decoupled.scala 218:16]
  reg  ram_last [0:15]; // @[Decoupled.scala 218:16]
  wire  ram_last_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16]
  wire [3:0] ram_last_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_last_MPORT_data; // @[Decoupled.scala 218:16]
  wire [3:0] ram_last_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_last_MPORT_mask; // @[Decoupled.scala 218:16]
  wire  ram_last_MPORT_en; // @[Decoupled.scala 218:16]
  reg [5:0] ram_mty [0:15]; // @[Decoupled.scala 218:16]
  wire [5:0] ram_mty_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16]
  wire [3:0] ram_mty_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16]
  wire [5:0] ram_mty_MPORT_data; // @[Decoupled.scala 218:16]
  wire [3:0] ram_mty_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_mty_MPORT_mask; // @[Decoupled.scala 218:16]
  wire  ram_mty_MPORT_en; // @[Decoupled.scala 218:16]
  reg [3:0] deq_ptr_value; // @[Counter.scala 60:40]
  wire  ptr_match = 4'h0 == deq_ptr_value; // @[Decoupled.scala 223:33]
  wire  do_deq = io_deq_ready & io_deq_valid; // @[Decoupled.scala 40:37]
  wire [3:0] _value_T_3 = deq_ptr_value + 4'h1; // @[Counter.scala 76:24]
  assign ram_data_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_data_io_deq_bits_MPORT_data = ram_data[ram_data_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  assign ram_data_MPORT_data = 512'h0;
  assign ram_data_MPORT_addr = 4'h0;
  assign ram_data_MPORT_mask = 1'h1;
  assign ram_data_MPORT_en = 1'h0;
  assign ram_tcrc_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_tcrc_io_deq_bits_MPORT_data = ram_tcrc[ram_tcrc_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  assign ram_tcrc_MPORT_data = 32'h0;
  assign ram_tcrc_MPORT_addr = 4'h0;
  assign ram_tcrc_MPORT_mask = 1'h1;
  assign ram_tcrc_MPORT_en = 1'h0;
  assign ram_ctrl_marker_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_ctrl_marker_io_deq_bits_MPORT_data = ram_ctrl_marker[ram_ctrl_marker_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  assign ram_ctrl_marker_MPORT_data = 1'h0;
  assign ram_ctrl_marker_MPORT_addr = 4'h0;
  assign ram_ctrl_marker_MPORT_mask = 1'h1;
  assign ram_ctrl_marker_MPORT_en = 1'h0;
  assign ram_ctrl_ecc_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_ctrl_ecc_io_deq_bits_MPORT_data = ram_ctrl_ecc[ram_ctrl_ecc_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  assign ram_ctrl_ecc_MPORT_data = 7'h0;
  assign ram_ctrl_ecc_MPORT_addr = 4'h0;
  assign ram_ctrl_ecc_MPORT_mask = 1'h1;
  assign ram_ctrl_ecc_MPORT_en = 1'h0;
  assign ram_ctrl_len_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_ctrl_len_io_deq_bits_MPORT_data = ram_ctrl_len[ram_ctrl_len_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  assign ram_ctrl_len_MPORT_data = 32'h0;
  assign ram_ctrl_len_MPORT_addr = 4'h0;
  assign ram_ctrl_len_MPORT_mask = 1'h1;
  assign ram_ctrl_len_MPORT_en = 1'h0;
  assign ram_ctrl_port_id_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_ctrl_port_id_io_deq_bits_MPORT_data = ram_ctrl_port_id[ram_ctrl_port_id_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  assign ram_ctrl_port_id_MPORT_data = 3'h0;
  assign ram_ctrl_port_id_MPORT_addr = 4'h0;
  assign ram_ctrl_port_id_MPORT_mask = 1'h1;
  assign ram_ctrl_port_id_MPORT_en = 1'h0;
  assign ram_ctrl_qid_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_ctrl_qid_io_deq_bits_MPORT_data = ram_ctrl_qid[ram_ctrl_qid_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  assign ram_ctrl_qid_MPORT_data = 11'h0;
  assign ram_ctrl_qid_MPORT_addr = 4'h0;
  assign ram_ctrl_qid_MPORT_mask = 1'h1;
  assign ram_ctrl_qid_MPORT_en = 1'h0;
  assign ram_ctrl_has_cmpt_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_ctrl_has_cmpt_io_deq_bits_MPORT_data = ram_ctrl_has_cmpt[ram_ctrl_has_cmpt_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  assign ram_ctrl_has_cmpt_MPORT_data = 1'h0;
  assign ram_ctrl_has_cmpt_MPORT_addr = 4'h0;
  assign ram_ctrl_has_cmpt_MPORT_mask = 1'h1;
  assign ram_ctrl_has_cmpt_MPORT_en = 1'h0;
  assign ram_last_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_last_io_deq_bits_MPORT_data = ram_last[ram_last_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  assign ram_last_MPORT_data = 1'h0;
  assign ram_last_MPORT_addr = 4'h0;
  assign ram_last_MPORT_mask = 1'h1;
  assign ram_last_MPORT_en = 1'h0;
  assign ram_mty_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_mty_io_deq_bits_MPORT_data = ram_mty[ram_mty_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  assign ram_mty_MPORT_data = 6'h0;
  assign ram_mty_MPORT_addr = 4'h0;
  assign ram_mty_MPORT_mask = 1'h1;
  assign ram_mty_MPORT_en = 1'h0;
  assign io_deq_valid = ~ptr_match; // @[Decoupled.scala 240:19]
  assign io_deq_bits_data = ram_data_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15]
  assign io_deq_bits_tcrc = ram_tcrc_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15]
  assign io_deq_bits_ctrl_marker = ram_ctrl_marker_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15]
  assign io_deq_bits_ctrl_ecc = ram_ctrl_ecc_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15]
  assign io_deq_bits_ctrl_len = ram_ctrl_len_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15]
  assign io_deq_bits_ctrl_port_id = ram_ctrl_port_id_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15]
  assign io_deq_bits_ctrl_qid = ram_ctrl_qid_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15]
  assign io_deq_bits_ctrl_has_cmpt = ram_ctrl_has_cmpt_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15]
  assign io_deq_bits_last = ram_last_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15]
  assign io_deq_bits_mty = ram_mty_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15]
  always @(posedge clock) begin
    if(ram_data_MPORT_en & ram_data_MPORT_mask) begin
      ram_data[ram_data_MPORT_addr] <= ram_data_MPORT_data; // @[Decoupled.scala 218:16]
    end
    if(ram_tcrc_MPORT_en & ram_tcrc_MPORT_mask) begin
      ram_tcrc[ram_tcrc_MPORT_addr] <= ram_tcrc_MPORT_data; // @[Decoupled.scala 218:16]
    end
    if(ram_ctrl_marker_MPORT_en & ram_ctrl_marker_MPORT_mask) begin
      ram_ctrl_marker[ram_ctrl_marker_MPORT_addr] <= ram_ctrl_marker_MPORT_data; // @[Decoupled.scala 218:16]
    end
    if(ram_ctrl_ecc_MPORT_en & ram_ctrl_ecc_MPORT_mask) begin
      ram_ctrl_ecc[ram_ctrl_ecc_MPORT_addr] <= ram_ctrl_ecc_MPORT_data; // @[Decoupled.scala 218:16]
    end
    if(ram_ctrl_len_MPORT_en & ram_ctrl_len_MPORT_mask) begin
      ram_ctrl_len[ram_ctrl_len_MPORT_addr] <= ram_ctrl_len_MPORT_data; // @[Decoupled.scala 218:16]
    end
    if(ram_ctrl_port_id_MPORT_en & ram_ctrl_port_id_MPORT_mask) begin
      ram_ctrl_port_id[ram_ctrl_port_id_MPORT_addr] <= ram_ctrl_port_id_MPORT_data; // @[Decoupled.scala 218:16]
    end
    if(ram_ctrl_qid_MPORT_en & ram_ctrl_qid_MPORT_mask) begin
      ram_ctrl_qid[ram_ctrl_qid_MPORT_addr] <= ram_ctrl_qid_MPORT_data; // @[Decoupled.scala 218:16]
    end
    if(ram_ctrl_has_cmpt_MPORT_en & ram_ctrl_has_cmpt_MPORT_mask) begin
      ram_ctrl_has_cmpt[ram_ctrl_has_cmpt_MPORT_addr] <= ram_ctrl_has_cmpt_MPORT_data; // @[Decoupled.scala 218:16]
    end
    if(ram_last_MPORT_en & ram_last_MPORT_mask) begin
      ram_last[ram_last_MPORT_addr] <= ram_last_MPORT_data; // @[Decoupled.scala 218:16]
    end
    if(ram_mty_MPORT_en & ram_mty_MPORT_mask) begin
      ram_mty[ram_mty_MPORT_addr] <= ram_mty_MPORT_data; // @[Decoupled.scala 218:16]
    end
    if (reset) begin // @[Counter.scala 60:40]
      deq_ptr_value <= 4'h0; // @[Counter.scala 60:40]
    end else if (do_deq) begin // @[Decoupled.scala 233:17]
      deq_ptr_value <= _value_T_3; // @[Counter.scala 76:15]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {16{`RANDOM}};
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    ram_data[initvar] = _RAND_0[511:0];
  _RAND_1 = {1{`RANDOM}};
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    ram_tcrc[initvar] = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    ram_ctrl_marker[initvar] = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    ram_ctrl_ecc[initvar] = _RAND_3[6:0];
  _RAND_4 = {1{`RANDOM}};
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    ram_ctrl_len[initvar] = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    ram_ctrl_port_id[initvar] = _RAND_5[2:0];
  _RAND_6 = {1{`RANDOM}};
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    ram_ctrl_qid[initvar] = _RAND_6[10:0];
  _RAND_7 = {1{`RANDOM}};
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    ram_ctrl_has_cmpt[initvar] = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    ram_last[initvar] = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    ram_mty[initvar] = _RAND_9[5:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  deq_ptr_value = _RAND_10[3:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module XQueue(
  input          clock,
  input          reset,
  input          io_out_ready,
  output         io_out_valid,
  output [511:0] io_out_bits_data,
  output [31:0]  io_out_bits_tcrc,
  output         io_out_bits_ctrl_marker,
  output [6:0]   io_out_bits_ctrl_ecc,
  output [31:0]  io_out_bits_ctrl_len,
  output [2:0]   io_out_bits_ctrl_port_id,
  output [10:0]  io_out_bits_ctrl_qid,
  output         io_out_bits_ctrl_has_cmpt,
  output         io_out_bits_last,
  output [5:0]   io_out_bits_mty
);
  wire  q_clock; // @[XQueue.scala 85:39]
  wire  q_reset; // @[XQueue.scala 85:39]
  wire  q_io_deq_ready; // @[XQueue.scala 85:39]
  wire  q_io_deq_valid; // @[XQueue.scala 85:39]
  wire [511:0] q_io_deq_bits_data; // @[XQueue.scala 85:39]
  wire [31:0] q_io_deq_bits_tcrc; // @[XQueue.scala 85:39]
  wire  q_io_deq_bits_ctrl_marker; // @[XQueue.scala 85:39]
  wire [6:0] q_io_deq_bits_ctrl_ecc; // @[XQueue.scala 85:39]
  wire [31:0] q_io_deq_bits_ctrl_len; // @[XQueue.scala 85:39]
  wire [2:0] q_io_deq_bits_ctrl_port_id; // @[XQueue.scala 85:39]
  wire [10:0] q_io_deq_bits_ctrl_qid; // @[XQueue.scala 85:39]
  wire  q_io_deq_bits_ctrl_has_cmpt; // @[XQueue.scala 85:39]
  wire  q_io_deq_bits_last; // @[XQueue.scala 85:39]
  wire [5:0] q_io_deq_bits_mty; // @[XQueue.scala 85:39]
  Queue_2 q ( // @[XQueue.scala 85:39]
    .clock(q_clock),
    .reset(q_reset),
    .io_deq_ready(q_io_deq_ready),
    .io_deq_valid(q_io_deq_valid),
    .io_deq_bits_data(q_io_deq_bits_data),
    .io_deq_bits_tcrc(q_io_deq_bits_tcrc),
    .io_deq_bits_ctrl_marker(q_io_deq_bits_ctrl_marker),
    .io_deq_bits_ctrl_ecc(q_io_deq_bits_ctrl_ecc),
    .io_deq_bits_ctrl_len(q_io_deq_bits_ctrl_len),
    .io_deq_bits_ctrl_port_id(q_io_deq_bits_ctrl_port_id),
    .io_deq_bits_ctrl_qid(q_io_deq_bits_ctrl_qid),
    .io_deq_bits_ctrl_has_cmpt(q_io_deq_bits_ctrl_has_cmpt),
    .io_deq_bits_last(q_io_deq_bits_last),
    .io_deq_bits_mty(q_io_deq_bits_mty)
  );
  assign io_out_valid = q_io_deq_valid; // @[XQueue.scala 88:34]
  assign io_out_bits_data = q_io_deq_bits_data; // @[XQueue.scala 88:34]
  assign io_out_bits_tcrc = q_io_deq_bits_tcrc; // @[XQueue.scala 88:34]
  assign io_out_bits_ctrl_marker = q_io_deq_bits_ctrl_marker; // @[XQueue.scala 88:34]
  assign io_out_bits_ctrl_ecc = q_io_deq_bits_ctrl_ecc; // @[XQueue.scala 88:34]
  assign io_out_bits_ctrl_len = q_io_deq_bits_ctrl_len; // @[XQueue.scala 88:34]
  assign io_out_bits_ctrl_port_id = q_io_deq_bits_ctrl_port_id; // @[XQueue.scala 88:34]
  assign io_out_bits_ctrl_qid = q_io_deq_bits_ctrl_qid; // @[XQueue.scala 88:34]
  assign io_out_bits_ctrl_has_cmpt = q_io_deq_bits_ctrl_has_cmpt; // @[XQueue.scala 88:34]
  assign io_out_bits_last = q_io_deq_bits_last; // @[XQueue.scala 88:34]
  assign io_out_bits_mty = q_io_deq_bits_mty; // @[XQueue.scala 88:34]
  assign q_clock = clock;
  assign q_reset = reset;
  assign q_io_deq_ready = io_out_ready; // @[XQueue.scala 88:34]
endmodule
module Queue_3(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input  [63:0] io_enq_bits_addr,
  input  [10:0] io_enq_bits_qid,
  input         io_enq_bits_error,
  input  [7:0]  io_enq_bits_func,
  input  [2:0]  io_enq_bits_port_id,
  input  [6:0]  io_enq_bits_pfch_tag,
  input  [31:0] io_enq_bits_len,
  input         io_deq_ready,
  output        io_deq_valid,
  output [63:0] io_deq_bits_addr,
  output [10:0] io_deq_bits_qid,
  output        io_deq_bits_error,
  output [7:0]  io_deq_bits_func,
  output [2:0]  io_deq_bits_port_id,
  output [6:0]  io_deq_bits_pfch_tag,
  output [31:0] io_deq_bits_len
);
`ifdef RANDOMIZE_MEM_INIT
  reg [63:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
`endif // RANDOMIZE_REG_INIT
  reg [63:0] ram_addr [0:15]; // @[Decoupled.scala 218:16]
  wire [63:0] ram_addr_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16]
  wire [3:0] ram_addr_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16]
  wire [63:0] ram_addr_MPORT_data; // @[Decoupled.scala 218:16]
  wire [3:0] ram_addr_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_addr_MPORT_mask; // @[Decoupled.scala 218:16]
  wire  ram_addr_MPORT_en; // @[Decoupled.scala 218:16]
  reg [10:0] ram_qid [0:15]; // @[Decoupled.scala 218:16]
  wire [10:0] ram_qid_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16]
  wire [3:0] ram_qid_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16]
  wire [10:0] ram_qid_MPORT_data; // @[Decoupled.scala 218:16]
  wire [3:0] ram_qid_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_qid_MPORT_mask; // @[Decoupled.scala 218:16]
  wire  ram_qid_MPORT_en; // @[Decoupled.scala 218:16]
  reg  ram_error [0:15]; // @[Decoupled.scala 218:16]
  wire  ram_error_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16]
  wire [3:0] ram_error_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_error_MPORT_data; // @[Decoupled.scala 218:16]
  wire [3:0] ram_error_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_error_MPORT_mask; // @[Decoupled.scala 218:16]
  wire  ram_error_MPORT_en; // @[Decoupled.scala 218:16]
  reg [7:0] ram_func [0:15]; // @[Decoupled.scala 218:16]
  wire [7:0] ram_func_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16]
  wire [3:0] ram_func_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16]
  wire [7:0] ram_func_MPORT_data; // @[Decoupled.scala 218:16]
  wire [3:0] ram_func_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_func_MPORT_mask; // @[Decoupled.scala 218:16]
  wire  ram_func_MPORT_en; // @[Decoupled.scala 218:16]
  reg [2:0] ram_port_id [0:15]; // @[Decoupled.scala 218:16]
  wire [2:0] ram_port_id_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16]
  wire [3:0] ram_port_id_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16]
  wire [2:0] ram_port_id_MPORT_data; // @[Decoupled.scala 218:16]
  wire [3:0] ram_port_id_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_port_id_MPORT_mask; // @[Decoupled.scala 218:16]
  wire  ram_port_id_MPORT_en; // @[Decoupled.scala 218:16]
  reg [6:0] ram_pfch_tag [0:15]; // @[Decoupled.scala 218:16]
  wire [6:0] ram_pfch_tag_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16]
  wire [3:0] ram_pfch_tag_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16]
  wire [6:0] ram_pfch_tag_MPORT_data; // @[Decoupled.scala 218:16]
  wire [3:0] ram_pfch_tag_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_pfch_tag_MPORT_mask; // @[Decoupled.scala 218:16]
  wire  ram_pfch_tag_MPORT_en; // @[Decoupled.scala 218:16]
  reg [31:0] ram_len [0:15]; // @[Decoupled.scala 218:16]
  wire [31:0] ram_len_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16]
  wire [3:0] ram_len_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16]
  wire [31:0] ram_len_MPORT_data; // @[Decoupled.scala 218:16]
  wire [3:0] ram_len_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_len_MPORT_mask; // @[Decoupled.scala 218:16]
  wire  ram_len_MPORT_en; // @[Decoupled.scala 218:16]
  reg [3:0] enq_ptr_value; // @[Counter.scala 60:40]
  reg [3:0] deq_ptr_value; // @[Counter.scala 60:40]
  reg  maybe_full; // @[Decoupled.scala 221:27]
  wire  ptr_match = enq_ptr_value == deq_ptr_value; // @[Decoupled.scala 223:33]
  wire  empty = ptr_match & ~maybe_full; // @[Decoupled.scala 224:25]
  wire  full = ptr_match & maybe_full; // @[Decoupled.scala 225:24]
  wire  do_enq = io_enq_ready & io_enq_valid; // @[Decoupled.scala 40:37]
  wire  do_deq = io_deq_ready & io_deq_valid; // @[Decoupled.scala 40:37]
  wire [3:0] _value_T_1 = enq_ptr_value + 4'h1; // @[Counter.scala 76:24]
  wire [3:0] _value_T_3 = deq_ptr_value + 4'h1; // @[Counter.scala 76:24]
  assign ram_addr_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_addr_io_deq_bits_MPORT_data = ram_addr[ram_addr_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  assign ram_addr_MPORT_data = io_enq_bits_addr;
  assign ram_addr_MPORT_addr = enq_ptr_value;
  assign ram_addr_MPORT_mask = 1'h1;
  assign ram_addr_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_qid_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_qid_io_deq_bits_MPORT_data = ram_qid[ram_qid_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  assign ram_qid_MPORT_data = io_enq_bits_qid;
  assign ram_qid_MPORT_addr = enq_ptr_value;
  assign ram_qid_MPORT_mask = 1'h1;
  assign ram_qid_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_error_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_error_io_deq_bits_MPORT_data = ram_error[ram_error_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  assign ram_error_MPORT_data = io_enq_bits_error;
  assign ram_error_MPORT_addr = enq_ptr_value;
  assign ram_error_MPORT_mask = 1'h1;
  assign ram_error_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_func_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_func_io_deq_bits_MPORT_data = ram_func[ram_func_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  assign ram_func_MPORT_data = io_enq_bits_func;
  assign ram_func_MPORT_addr = enq_ptr_value;
  assign ram_func_MPORT_mask = 1'h1;
  assign ram_func_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_port_id_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_port_id_io_deq_bits_MPORT_data = ram_port_id[ram_port_id_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  assign ram_port_id_MPORT_data = io_enq_bits_port_id;
  assign ram_port_id_MPORT_addr = enq_ptr_value;
  assign ram_port_id_MPORT_mask = 1'h1;
  assign ram_port_id_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_pfch_tag_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_pfch_tag_io_deq_bits_MPORT_data = ram_pfch_tag[ram_pfch_tag_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  assign ram_pfch_tag_MPORT_data = io_enq_bits_pfch_tag;
  assign ram_pfch_tag_MPORT_addr = enq_ptr_value;
  assign ram_pfch_tag_MPORT_mask = 1'h1;
  assign ram_pfch_tag_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_len_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_len_io_deq_bits_MPORT_data = ram_len[ram_len_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  assign ram_len_MPORT_data = io_enq_bits_len;
  assign ram_len_MPORT_addr = enq_ptr_value;
  assign ram_len_MPORT_mask = 1'h1;
  assign ram_len_MPORT_en = io_enq_ready & io_enq_valid;
  assign io_enq_ready = ~full; // @[Decoupled.scala 241:19]
  assign io_deq_valid = ~empty; // @[Decoupled.scala 240:19]
  assign io_deq_bits_addr = ram_addr_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15]
  assign io_deq_bits_qid = ram_qid_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15]
  assign io_deq_bits_error = ram_error_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15]
  assign io_deq_bits_func = ram_func_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15]
  assign io_deq_bits_port_id = ram_port_id_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15]
  assign io_deq_bits_pfch_tag = ram_pfch_tag_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15]
  assign io_deq_bits_len = ram_len_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15]
  always @(posedge clock) begin
    if(ram_addr_MPORT_en & ram_addr_MPORT_mask) begin
      ram_addr[ram_addr_MPORT_addr] <= ram_addr_MPORT_data; // @[Decoupled.scala 218:16]
    end
    if(ram_qid_MPORT_en & ram_qid_MPORT_mask) begin
      ram_qid[ram_qid_MPORT_addr] <= ram_qid_MPORT_data; // @[Decoupled.scala 218:16]
    end
    if(ram_error_MPORT_en & ram_error_MPORT_mask) begin
      ram_error[ram_error_MPORT_addr] <= ram_error_MPORT_data; // @[Decoupled.scala 218:16]
    end
    if(ram_func_MPORT_en & ram_func_MPORT_mask) begin
      ram_func[ram_func_MPORT_addr] <= ram_func_MPORT_data; // @[Decoupled.scala 218:16]
    end
    if(ram_port_id_MPORT_en & ram_port_id_MPORT_mask) begin
      ram_port_id[ram_port_id_MPORT_addr] <= ram_port_id_MPORT_data; // @[Decoupled.scala 218:16]
    end
    if(ram_pfch_tag_MPORT_en & ram_pfch_tag_MPORT_mask) begin
      ram_pfch_tag[ram_pfch_tag_MPORT_addr] <= ram_pfch_tag_MPORT_data; // @[Decoupled.scala 218:16]
    end
    if(ram_len_MPORT_en & ram_len_MPORT_mask) begin
      ram_len[ram_len_MPORT_addr] <= ram_len_MPORT_data; // @[Decoupled.scala 218:16]
    end
    if (reset) begin // @[Counter.scala 60:40]
      enq_ptr_value <= 4'h0; // @[Counter.scala 60:40]
    end else if (do_enq) begin // @[Decoupled.scala 229:17]
      enq_ptr_value <= _value_T_1; // @[Counter.scala 76:15]
    end
    if (reset) begin // @[Counter.scala 60:40]
      deq_ptr_value <= 4'h0; // @[Counter.scala 60:40]
    end else if (do_deq) begin // @[Decoupled.scala 233:17]
      deq_ptr_value <= _value_T_3; // @[Counter.scala 76:15]
    end
    if (reset) begin // @[Decoupled.scala 221:27]
      maybe_full <= 1'h0; // @[Decoupled.scala 221:27]
    end else if (do_enq != do_deq) begin // @[Decoupled.scala 236:28]
      maybe_full <= do_enq; // @[Decoupled.scala 237:16]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {2{`RANDOM}};
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    ram_addr[initvar] = _RAND_0[63:0];
  _RAND_1 = {1{`RANDOM}};
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    ram_qid[initvar] = _RAND_1[10:0];
  _RAND_2 = {1{`RANDOM}};
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    ram_error[initvar] = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    ram_func[initvar] = _RAND_3[7:0];
  _RAND_4 = {1{`RANDOM}};
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    ram_port_id[initvar] = _RAND_4[2:0];
  _RAND_5 = {1{`RANDOM}};
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    ram_pfch_tag[initvar] = _RAND_5[6:0];
  _RAND_6 = {1{`RANDOM}};
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    ram_len[initvar] = _RAND_6[31:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  enq_ptr_value = _RAND_7[3:0];
  _RAND_8 = {1{`RANDOM}};
  deq_ptr_value = _RAND_8[3:0];
  _RAND_9 = {1{`RANDOM}};
  maybe_full = _RAND_9[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module XQueue_1(
  input         clock,
  input         reset,
  output        io_in_ready,
  input         io_in_valid,
  input  [63:0] io_in_bits_addr,
  input  [10:0] io_in_bits_qid,
  input         io_in_bits_error,
  input  [7:0]  io_in_bits_func,
  input  [2:0]  io_in_bits_port_id,
  input  [6:0]  io_in_bits_pfch_tag,
  input  [31:0] io_in_bits_len,
  input         io_out_ready,
  output        io_out_valid,
  output [63:0] io_out_bits_addr,
  output [10:0] io_out_bits_qid,
  output        io_out_bits_error,
  output [7:0]  io_out_bits_func,
  output [2:0]  io_out_bits_port_id,
  output [6:0]  io_out_bits_pfch_tag,
  output [31:0] io_out_bits_len
);
  wire  q_clock; // @[XQueue.scala 85:39]
  wire  q_reset; // @[XQueue.scala 85:39]
  wire  q_io_enq_ready; // @[XQueue.scala 85:39]
  wire  q_io_enq_valid; // @[XQueue.scala 85:39]
  wire [63:0] q_io_enq_bits_addr; // @[XQueue.scala 85:39]
  wire [10:0] q_io_enq_bits_qid; // @[XQueue.scala 85:39]
  wire  q_io_enq_bits_error; // @[XQueue.scala 85:39]
  wire [7:0] q_io_enq_bits_func; // @[XQueue.scala 85:39]
  wire [2:0] q_io_enq_bits_port_id; // @[XQueue.scala 85:39]
  wire [6:0] q_io_enq_bits_pfch_tag; // @[XQueue.scala 85:39]
  wire [31:0] q_io_enq_bits_len; // @[XQueue.scala 85:39]
  wire  q_io_deq_ready; // @[XQueue.scala 85:39]
  wire  q_io_deq_valid; // @[XQueue.scala 85:39]
  wire [63:0] q_io_deq_bits_addr; // @[XQueue.scala 85:39]
  wire [10:0] q_io_deq_bits_qid; // @[XQueue.scala 85:39]
  wire  q_io_deq_bits_error; // @[XQueue.scala 85:39]
  wire [7:0] q_io_deq_bits_func; // @[XQueue.scala 85:39]
  wire [2:0] q_io_deq_bits_port_id; // @[XQueue.scala 85:39]
  wire [6:0] q_io_deq_bits_pfch_tag; // @[XQueue.scala 85:39]
  wire [31:0] q_io_deq_bits_len; // @[XQueue.scala 85:39]
  Queue_3 q ( // @[XQueue.scala 85:39]
    .clock(q_clock),
    .reset(q_reset),
    .io_enq_ready(q_io_enq_ready),
    .io_enq_valid(q_io_enq_valid),
    .io_enq_bits_addr(q_io_enq_bits_addr),
    .io_enq_bits_qid(q_io_enq_bits_qid),
    .io_enq_bits_error(q_io_enq_bits_error),
    .io_enq_bits_func(q_io_enq_bits_func),
    .io_enq_bits_port_id(q_io_enq_bits_port_id),
    .io_enq_bits_pfch_tag(q_io_enq_bits_pfch_tag),
    .io_enq_bits_len(q_io_enq_bits_len),
    .io_deq_ready(q_io_deq_ready),
    .io_deq_valid(q_io_deq_valid),
    .io_deq_bits_addr(q_io_deq_bits_addr),
    .io_deq_bits_qid(q_io_deq_bits_qid),
    .io_deq_bits_error(q_io_deq_bits_error),
    .io_deq_bits_func(q_io_deq_bits_func),
    .io_deq_bits_port_id(q_io_deq_bits_port_id),
    .io_deq_bits_pfch_tag(q_io_deq_bits_pfch_tag),
    .io_deq_bits_len(q_io_deq_bits_len)
  );
  assign io_in_ready = q_io_enq_ready; // @[XQueue.scala 87:34]
  assign io_out_valid = q_io_deq_valid; // @[XQueue.scala 88:34]
  assign io_out_bits_addr = q_io_deq_bits_addr; // @[XQueue.scala 88:34]
  assign io_out_bits_qid = q_io_deq_bits_qid; // @[XQueue.scala 88:34]
  assign io_out_bits_error = q_io_deq_bits_error; // @[XQueue.scala 88:34]
  assign io_out_bits_func = q_io_deq_bits_func; // @[XQueue.scala 88:34]
  assign io_out_bits_port_id = q_io_deq_bits_port_id; // @[XQueue.scala 88:34]
  assign io_out_bits_pfch_tag = q_io_deq_bits_pfch_tag; // @[XQueue.scala 88:34]
  assign io_out_bits_len = q_io_deq_bits_len; // @[XQueue.scala 88:34]
  assign q_clock = clock;
  assign q_reset = reset;
  assign q_io_enq_valid = io_in_valid; // @[XQueue.scala 87:34]
  assign q_io_enq_bits_addr = io_in_bits_addr; // @[XQueue.scala 87:34]
  assign q_io_enq_bits_qid = io_in_bits_qid; // @[XQueue.scala 87:34]
  assign q_io_enq_bits_error = io_in_bits_error; // @[XQueue.scala 87:34]
  assign q_io_enq_bits_func = io_in_bits_func; // @[XQueue.scala 87:34]
  assign q_io_enq_bits_port_id = io_in_bits_port_id; // @[XQueue.scala 87:34]
  assign q_io_enq_bits_pfch_tag = io_in_bits_pfch_tag; // @[XQueue.scala 87:34]
  assign q_io_enq_bits_len = io_in_bits_len; // @[XQueue.scala 87:34]
  assign q_io_deq_ready = io_out_ready; // @[XQueue.scala 88:34]
endmodule
module DataBoundarySplit(
  input          clock,
  input          reset,
  output         io_cmd_in_ready,
  input          io_cmd_in_valid,
  input  [63:0]  io_cmd_in_bits_addr,
  input  [10:0]  io_cmd_in_bits_qid,
  input          io_cmd_in_bits_error,
  input  [7:0]   io_cmd_in_bits_func,
  input  [2:0]   io_cmd_in_bits_port_id,
  input  [6:0]   io_cmd_in_bits_pfch_tag,
  input  [31:0]  io_cmd_in_bits_len,
  input          io_data_out_ready,
  output         io_data_out_valid,
  output [511:0] io_data_out_bits_data,
  output [31:0]  io_data_out_bits_tcrc,
  output         io_data_out_bits_ctrl_marker,
  output [6:0]   io_data_out_bits_ctrl_ecc,
  output [31:0]  io_data_out_bits_ctrl_len,
  output [2:0]   io_data_out_bits_ctrl_port_id,
  output [10:0]  io_data_out_bits_ctrl_qid,
  output         io_data_out_bits_ctrl_has_cmpt,
  output         io_data_out_bits_last,
  output [5:0]   io_data_out_bits_mty,
  input          io_cmd_out_ready,
  output         io_cmd_out_valid,
  output [63:0]  io_cmd_out_bits_addr,
  output [10:0]  io_cmd_out_bits_qid,
  output         io_cmd_out_bits_error,
  output [7:0]   io_cmd_out_bits_func,
  output [2:0]   io_cmd_out_bits_port_id,
  output [6:0]   io_cmd_out_bits_pfch_tag,
  output [31:0]  io_cmd_out_bits_len
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire  data_fifo_clock; // @[XQueue.scala 35:23]
  wire  data_fifo_reset; // @[XQueue.scala 35:23]
  wire  data_fifo_io_out_ready; // @[XQueue.scala 35:23]
  wire  data_fifo_io_out_valid; // @[XQueue.scala 35:23]
  wire [511:0] data_fifo_io_out_bits_data; // @[XQueue.scala 35:23]
  wire [31:0] data_fifo_io_out_bits_tcrc; // @[XQueue.scala 35:23]
  wire  data_fifo_io_out_bits_ctrl_marker; // @[XQueue.scala 35:23]
  wire [6:0] data_fifo_io_out_bits_ctrl_ecc; // @[XQueue.scala 35:23]
  wire [31:0] data_fifo_io_out_bits_ctrl_len; // @[XQueue.scala 35:23]
  wire [2:0] data_fifo_io_out_bits_ctrl_port_id; // @[XQueue.scala 35:23]
  wire [10:0] data_fifo_io_out_bits_ctrl_qid; // @[XQueue.scala 35:23]
  wire  data_fifo_io_out_bits_ctrl_has_cmpt; // @[XQueue.scala 35:23]
  wire  data_fifo_io_out_bits_last; // @[XQueue.scala 35:23]
  wire [5:0] data_fifo_io_out_bits_mty; // @[XQueue.scala 35:23]
  wire  cmd_fifo_clock; // @[XQueue.scala 35:23]
  wire  cmd_fifo_reset; // @[XQueue.scala 35:23]
  wire  cmd_fifo_io_in_ready; // @[XQueue.scala 35:23]
  wire  cmd_fifo_io_in_valid; // @[XQueue.scala 35:23]
  wire [63:0] cmd_fifo_io_in_bits_addr; // @[XQueue.scala 35:23]
  wire [10:0] cmd_fifo_io_in_bits_qid; // @[XQueue.scala 35:23]
  wire  cmd_fifo_io_in_bits_error; // @[XQueue.scala 35:23]
  wire [7:0] cmd_fifo_io_in_bits_func; // @[XQueue.scala 35:23]
  wire [2:0] cmd_fifo_io_in_bits_port_id; // @[XQueue.scala 35:23]
  wire [6:0] cmd_fifo_io_in_bits_pfch_tag; // @[XQueue.scala 35:23]
  wire [31:0] cmd_fifo_io_in_bits_len; // @[XQueue.scala 35:23]
  wire  cmd_fifo_io_out_ready; // @[XQueue.scala 35:23]
  wire  cmd_fifo_io_out_valid; // @[XQueue.scala 35:23]
  wire [63:0] cmd_fifo_io_out_bits_addr; // @[XQueue.scala 35:23]
  wire [10:0] cmd_fifo_io_out_bits_qid; // @[XQueue.scala 35:23]
  wire  cmd_fifo_io_out_bits_error; // @[XQueue.scala 35:23]
  wire [7:0] cmd_fifo_io_out_bits_func; // @[XQueue.scala 35:23]
  wire [2:0] cmd_fifo_io_out_bits_port_id; // @[XQueue.scala 35:23]
  wire [6:0] cmd_fifo_io_out_bits_pfch_tag; // @[XQueue.scala 35:23]
  wire [31:0] cmd_fifo_io_out_bits_len; // @[XQueue.scala 35:23]
  reg  state; // @[CheckSplit.scala 27:50]
  wire  _io_cmd_in_ready_T = ~state; // @[CheckSplit.scala 29:67]
  wire  _T_1 = io_cmd_in_ready & io_cmd_in_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_7 = _T_1 | state; // @[CheckSplit.scala 39:47 CheckSplit.scala 41:41 CheckSplit.scala 27:50]
  wire [31:0] _GEN_9 = _T_1 ? io_cmd_in_bits_len : 32'h0; // @[CheckSplit.scala 39:47 CheckSplit.scala 43:65 CheckSplit.scala 35:65]
  wire [6:0] _GEN_10 = _T_1 ? io_cmd_in_bits_pfch_tag : 7'h0; // @[CheckSplit.scala 39:47 CheckSplit.scala 43:65 CheckSplit.scala 35:65]
  wire [2:0] _GEN_11 = _T_1 ? io_cmd_in_bits_port_id : 3'h0; // @[CheckSplit.scala 39:47 CheckSplit.scala 43:65 CheckSplit.scala 35:65]
  wire [7:0] _GEN_12 = _T_1 ? io_cmd_in_bits_func : 8'h0; // @[CheckSplit.scala 39:47 CheckSplit.scala 43:65 CheckSplit.scala 35:65]
  wire  _GEN_13 = _T_1 & io_cmd_in_bits_error; // @[CheckSplit.scala 39:47 CheckSplit.scala 43:65 CheckSplit.scala 35:65]
  wire [10:0] _GEN_14 = _T_1 ? io_cmd_in_bits_qid : 11'h0; // @[CheckSplit.scala 39:47 CheckSplit.scala 43:65 CheckSplit.scala 35:65]
  wire [63:0] _GEN_15 = _T_1 ? io_cmd_in_bits_addr : 64'h0; // @[CheckSplit.scala 39:47 CheckSplit.scala 43:65 CheckSplit.scala 35:65]
  XQueue data_fifo ( // @[XQueue.scala 35:23]
    .clock(data_fifo_clock),
    .reset(data_fifo_reset),
    .io_out_ready(data_fifo_io_out_ready),
    .io_out_valid(data_fifo_io_out_valid),
    .io_out_bits_data(data_fifo_io_out_bits_data),
    .io_out_bits_tcrc(data_fifo_io_out_bits_tcrc),
    .io_out_bits_ctrl_marker(data_fifo_io_out_bits_ctrl_marker),
    .io_out_bits_ctrl_ecc(data_fifo_io_out_bits_ctrl_ecc),
    .io_out_bits_ctrl_len(data_fifo_io_out_bits_ctrl_len),
    .io_out_bits_ctrl_port_id(data_fifo_io_out_bits_ctrl_port_id),
    .io_out_bits_ctrl_qid(data_fifo_io_out_bits_ctrl_qid),
    .io_out_bits_ctrl_has_cmpt(data_fifo_io_out_bits_ctrl_has_cmpt),
    .io_out_bits_last(data_fifo_io_out_bits_last),
    .io_out_bits_mty(data_fifo_io_out_bits_mty)
  );
  XQueue_1 cmd_fifo ( // @[XQueue.scala 35:23]
    .clock(cmd_fifo_clock),
    .reset(cmd_fifo_reset),
    .io_in_ready(cmd_fifo_io_in_ready),
    .io_in_valid(cmd_fifo_io_in_valid),
    .io_in_bits_addr(cmd_fifo_io_in_bits_addr),
    .io_in_bits_qid(cmd_fifo_io_in_bits_qid),
    .io_in_bits_error(cmd_fifo_io_in_bits_error),
    .io_in_bits_func(cmd_fifo_io_in_bits_func),
    .io_in_bits_port_id(cmd_fifo_io_in_bits_port_id),
    .io_in_bits_pfch_tag(cmd_fifo_io_in_bits_pfch_tag),
    .io_in_bits_len(cmd_fifo_io_in_bits_len),
    .io_out_ready(cmd_fifo_io_out_ready),
    .io_out_valid(cmd_fifo_io_out_valid),
    .io_out_bits_addr(cmd_fifo_io_out_bits_addr),
    .io_out_bits_qid(cmd_fifo_io_out_bits_qid),
    .io_out_bits_error(cmd_fifo_io_out_bits_error),
    .io_out_bits_func(cmd_fifo_io_out_bits_func),
    .io_out_bits_port_id(cmd_fifo_io_out_bits_port_id),
    .io_out_bits_pfch_tag(cmd_fifo_io_out_bits_pfch_tag),
    .io_out_bits_len(cmd_fifo_io_out_bits_len)
  );
  assign io_cmd_in_ready = ~state & cmd_fifo_io_in_ready; // @[CheckSplit.scala 29:78]
  assign io_data_out_valid = data_fifo_io_out_valid; // @[CheckSplit.scala 23:25]
  assign io_data_out_bits_data = data_fifo_io_out_bits_data; // @[CheckSplit.scala 23:25]
  assign io_data_out_bits_tcrc = data_fifo_io_out_bits_tcrc; // @[CheckSplit.scala 23:25]
  assign io_data_out_bits_ctrl_marker = data_fifo_io_out_bits_ctrl_marker; // @[CheckSplit.scala 23:25]
  assign io_data_out_bits_ctrl_ecc = data_fifo_io_out_bits_ctrl_ecc; // @[CheckSplit.scala 23:25]
  assign io_data_out_bits_ctrl_len = data_fifo_io_out_bits_ctrl_len; // @[CheckSplit.scala 23:25]
  assign io_data_out_bits_ctrl_port_id = data_fifo_io_out_bits_ctrl_port_id; // @[CheckSplit.scala 23:25]
  assign io_data_out_bits_ctrl_qid = data_fifo_io_out_bits_ctrl_qid; // @[CheckSplit.scala 23:25]
  assign io_data_out_bits_ctrl_has_cmpt = data_fifo_io_out_bits_ctrl_has_cmpt; // @[CheckSplit.scala 23:25]
  assign io_data_out_bits_last = data_fifo_io_out_bits_last; // @[CheckSplit.scala 23:25]
  assign io_data_out_bits_mty = data_fifo_io_out_bits_mty; // @[CheckSplit.scala 23:25]
  assign io_cmd_out_valid = cmd_fifo_io_out_valid; // @[CheckSplit.scala 24:25]
  assign io_cmd_out_bits_addr = cmd_fifo_io_out_bits_addr; // @[CheckSplit.scala 24:25]
  assign io_cmd_out_bits_qid = cmd_fifo_io_out_bits_qid; // @[CheckSplit.scala 24:25]
  assign io_cmd_out_bits_error = cmd_fifo_io_out_bits_error; // @[CheckSplit.scala 24:25]
  assign io_cmd_out_bits_func = cmd_fifo_io_out_bits_func; // @[CheckSplit.scala 24:25]
  assign io_cmd_out_bits_port_id = cmd_fifo_io_out_bits_port_id; // @[CheckSplit.scala 24:25]
  assign io_cmd_out_bits_pfch_tag = cmd_fifo_io_out_bits_pfch_tag; // @[CheckSplit.scala 24:25]
  assign io_cmd_out_bits_len = cmd_fifo_io_out_bits_len; // @[CheckSplit.scala 24:25]
  assign data_fifo_clock = clock;
  assign data_fifo_reset = reset;
  assign data_fifo_io_out_ready = io_data_out_ready; // @[CheckSplit.scala 23:25]
  assign cmd_fifo_clock = clock;
  assign cmd_fifo_reset = reset;
  assign cmd_fifo_io_in_valid = _io_cmd_in_ready_T & _T_1; // @[Conditional.scala 40:58 CheckSplit.scala 34:57]
  assign cmd_fifo_io_in_bits_addr = _io_cmd_in_ready_T ? _GEN_15 : 64'h0; // @[Conditional.scala 40:58 CheckSplit.scala 35:65]
  assign cmd_fifo_io_in_bits_qid = _io_cmd_in_ready_T ? _GEN_14 : 11'h0; // @[Conditional.scala 40:58 CheckSplit.scala 35:65]
  assign cmd_fifo_io_in_bits_error = _io_cmd_in_ready_T & _GEN_13; // @[Conditional.scala 40:58 CheckSplit.scala 35:65]
  assign cmd_fifo_io_in_bits_func = _io_cmd_in_ready_T ? _GEN_12 : 8'h0; // @[Conditional.scala 40:58 CheckSplit.scala 35:65]
  assign cmd_fifo_io_in_bits_port_id = _io_cmd_in_ready_T ? _GEN_11 : 3'h0; // @[Conditional.scala 40:58 CheckSplit.scala 35:65]
  assign cmd_fifo_io_in_bits_pfch_tag = _io_cmd_in_ready_T ? _GEN_10 : 7'h0; // @[Conditional.scala 40:58 CheckSplit.scala 35:65]
  assign cmd_fifo_io_in_bits_len = _io_cmd_in_ready_T ? _GEN_9 : 32'h0; // @[Conditional.scala 40:58 CheckSplit.scala 35:65]
  assign cmd_fifo_io_out_ready = io_cmd_out_ready; // @[CheckSplit.scala 24:25]
  always @(posedge clock) begin
    if (reset) begin // @[CheckSplit.scala 27:50]
      state <= 1'h0; // @[CheckSplit.scala 27:50]
    end else if (_io_cmd_in_ready_T) begin // @[Conditional.scala 40:58]
      state <= _GEN_7;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module QDMADynamic(
  input          io_qdma_port_axi_aclk,
  input          io_qdma_port_axi_aresetn,
  input  [3:0]   io_qdma_port_m_axib_awid,
  input  [63:0]  io_qdma_port_m_axib_awaddr,
  input  [7:0]   io_qdma_port_m_axib_awlen,
  input  [2:0]   io_qdma_port_m_axib_awsize,
  input  [1:0]   io_qdma_port_m_axib_awburst,
  input  [2:0]   io_qdma_port_m_axib_awprot,
  input          io_qdma_port_m_axib_awlock,
  input  [3:0]   io_qdma_port_m_axib_awcache,
  input          io_qdma_port_m_axib_awvalid,
  output         io_qdma_port_m_axib_awready,
  input  [511:0] io_qdma_port_m_axib_wdata,
  input  [63:0]  io_qdma_port_m_axib_wstrb,
  input          io_qdma_port_m_axib_wlast,
  input          io_qdma_port_m_axib_wvalid,
  output         io_qdma_port_m_axib_wready,
  output [3:0]   io_qdma_port_m_axib_bid,
  output [1:0]   io_qdma_port_m_axib_bresp,
  output         io_qdma_port_m_axib_bvalid,
  input          io_qdma_port_m_axib_bready,
  input  [3:0]   io_qdma_port_m_axib_arid,
  input  [63:0]  io_qdma_port_m_axib_araddr,
  input  [7:0]   io_qdma_port_m_axib_arlen,
  input  [2:0]   io_qdma_port_m_axib_arsize,
  input  [1:0]   io_qdma_port_m_axib_arburst,
  input  [2:0]   io_qdma_port_m_axib_arprot,
  input          io_qdma_port_m_axib_arlock,
  input  [3:0]   io_qdma_port_m_axib_arcache,
  input          io_qdma_port_m_axib_arvalid,
  output         io_qdma_port_m_axib_arready,
  output [3:0]   io_qdma_port_m_axib_rid,
  output [511:0] io_qdma_port_m_axib_rdata,
  output [1:0]   io_qdma_port_m_axib_rresp,
  output         io_qdma_port_m_axib_rlast,
  output         io_qdma_port_m_axib_rvalid,
  input          io_qdma_port_m_axib_rready,
  input  [31:0]  io_qdma_port_m_axil_awaddr,
  input          io_qdma_port_m_axil_awvalid,
  output         io_qdma_port_m_axil_awready,
  input  [31:0]  io_qdma_port_m_axil_wdata,
  input  [3:0]   io_qdma_port_m_axil_wstrb,
  input          io_qdma_port_m_axil_wvalid,
  output         io_qdma_port_m_axil_wready,
  output [1:0]   io_qdma_port_m_axil_bresp,
  output         io_qdma_port_m_axil_bvalid,
  input          io_qdma_port_m_axil_bready,
  input  [31:0]  io_qdma_port_m_axil_araddr,
  input          io_qdma_port_m_axil_arvalid,
  output         io_qdma_port_m_axil_arready,
  output [31:0]  io_qdma_port_m_axil_rdata,
  output [1:0]   io_qdma_port_m_axil_rresp,
  output         io_qdma_port_m_axil_rvalid,
  input          io_qdma_port_m_axil_rready,
  output [63:0]  io_qdma_port_h2c_byp_in_st_addr,
  output [31:0]  io_qdma_port_h2c_byp_in_st_len,
  output         io_qdma_port_h2c_byp_in_st_eop,
  output         io_qdma_port_h2c_byp_in_st_sop,
  output         io_qdma_port_h2c_byp_in_st_mrkr_req,
  output         io_qdma_port_h2c_byp_in_st_sdi,
  output [10:0]  io_qdma_port_h2c_byp_in_st_qid,
  output         io_qdma_port_h2c_byp_in_st_error,
  output [7:0]   io_qdma_port_h2c_byp_in_st_func,
  output [15:0]  io_qdma_port_h2c_byp_in_st_cidx,
  output [2:0]   io_qdma_port_h2c_byp_in_st_port_id,
  output         io_qdma_port_h2c_byp_in_st_no_dma,
  output         io_qdma_port_h2c_byp_in_st_vld,
  input          io_qdma_port_h2c_byp_in_st_rdy,
  output [63:0]  io_qdma_port_c2h_byp_in_st_csh_addr,
  output [10:0]  io_qdma_port_c2h_byp_in_st_csh_qid,
  output         io_qdma_port_c2h_byp_in_st_csh_error,
  output [7:0]   io_qdma_port_c2h_byp_in_st_csh_func,
  output [2:0]   io_qdma_port_c2h_byp_in_st_csh_port_id,
  output [6:0]   io_qdma_port_c2h_byp_in_st_csh_pfch_tag,
  output         io_qdma_port_c2h_byp_in_st_csh_vld,
  input          io_qdma_port_c2h_byp_in_st_csh_rdy,
  output [511:0] io_qdma_port_s_axis_c2h_tdata,
  output [31:0]  io_qdma_port_s_axis_c2h_tcrc,
  output         io_qdma_port_s_axis_c2h_ctrl_marker,
  output [6:0]   io_qdma_port_s_axis_c2h_ctrl_ecc,
  output [31:0]  io_qdma_port_s_axis_c2h_ctrl_len,
  output [2:0]   io_qdma_port_s_axis_c2h_ctrl_port_id,
  output [10:0]  io_qdma_port_s_axis_c2h_ctrl_qid,
  output         io_qdma_port_s_axis_c2h_ctrl_has_cmpt,
  output [5:0]   io_qdma_port_s_axis_c2h_mty,
  output         io_qdma_port_s_axis_c2h_tlast,
  output         io_qdma_port_s_axis_c2h_tvalid,
  input          io_qdma_port_s_axis_c2h_tready,
  input  [511:0] io_qdma_port_m_axis_h2c_tdata,
  input  [31:0]  io_qdma_port_m_axis_h2c_tcrc,
  input  [10:0]  io_qdma_port_m_axis_h2c_tuser_qid,
  input  [2:0]   io_qdma_port_m_axis_h2c_tuser_port_id,
  input          io_qdma_port_m_axis_h2c_tuser_err,
  input  [31:0]  io_qdma_port_m_axis_h2c_tuser_mdata,
  input  [5:0]   io_qdma_port_m_axis_h2c_tuser_mty,
  input          io_qdma_port_m_axis_h2c_tuser_zero_byte,
  input          io_qdma_port_m_axis_h2c_tlast,
  input          io_qdma_port_m_axis_h2c_tvalid,
  output         io_qdma_port_m_axis_h2c_tready,
  input          io_user_clk,
  input          io_user_arstn,
  output         io_h2c_cmd_ready,
  input          io_h2c_cmd_valid,
  input  [63:0]  io_h2c_cmd_bits_addr,
  input  [31:0]  io_h2c_cmd_bits_len,
  output         io_h2c_data_valid,
  output [31:0]  io_reg_control_0,
  output [31:0]  io_reg_control_8,
  output [31:0]  io_reg_control_9,
  output [31:0]  io_reg_control_10,
  output [31:0]  io_reg_control_11,
  output [31:0]  io_reg_control_12,
  output [31:0]  io_reg_control_13,
  output [31:0]  io_reg_control_14,
  input  [31:0]  io_reg_status_300,
  input  [31:0]  io_reg_status_400,
  input  [31:0]  io_reg_status_401,
  input  [31:0]  io_reg_status_402,
  input  [31:0]  io_reg_status_403,
  input  [31:0]  io_reg_status_404,
  input  [31:0]  io_reg_status_405,
  input  [31:0]  io_reg_status_406,
  input  [31:0]  io_reg_status_407,
  input  [31:0]  io_reg_status_408,
  input  [31:0]  io_reg_status_409,
  input  [31:0]  io_reg_status_410,
  input  [31:0]  io_reg_status_411,
  input  [31:0]  io_reg_status_412,
  input  [31:0]  io_reg_status_413,
  input  [31:0]  io_reg_status_414,
  input          io_axib_aw_ready,
  output         io_axib_aw_valid,
  output [63:0]  io_axib_aw_bits_addr,
  input          io_axib_w_ready,
  output         io_axib_w_valid,
  output [511:0] io_axib_w_bits_data,
  output         io_axib_r_ready,
  input  [511:0] io_axib_r_bits_data,
  output         io_out_valid,
  output [31:0]  counter_4_0,
  output         io_out_ready,
  output [31:0]  counter_7_0,
  output [31:0]  counter_1_0,
  output         io_in_ready,
  output [31:0]  counter_3_1,
  output         io_out_ready_0,
  output [31:0]  counter_6_0,
  output         io_out_valid_0,
  output [31:0]  counter_0,
  output         io_in_valid,
  output [31:0]  io_tlb_miss_count,
  output         io_out_valid_1,
  output [31:0]  counter_2_1,
  output [31:0]  counter_5_0,
  output         io_out_ready_1
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
`endif // RANDOMIZE_REG_INIT
  wire  sw_reset_pad_O; // @[Buf.scala 33:34]
  wire  sw_reset_pad_I; // @[Buf.scala 33:34]
  wire  fifo_h2c_data_io__in_clk; // @[XConverter.scala 61:33]
  wire  fifo_h2c_data_io__out_clk; // @[XConverter.scala 61:33]
  wire  fifo_h2c_data_io__rstn; // @[XConverter.scala 61:33]
  wire  fifo_h2c_data_io__in_ready; // @[XConverter.scala 61:33]
  wire  fifo_h2c_data_io__in_valid; // @[XConverter.scala 61:33]
  wire [511:0] fifo_h2c_data_io__in_bits_data; // @[XConverter.scala 61:33]
  wire [31:0] fifo_h2c_data_io__in_bits_tcrc; // @[XConverter.scala 61:33]
  wire [10:0] fifo_h2c_data_io__in_bits_tuser_qid; // @[XConverter.scala 61:33]
  wire [2:0] fifo_h2c_data_io__in_bits_tuser_port_id; // @[XConverter.scala 61:33]
  wire  fifo_h2c_data_io__in_bits_tuser_err; // @[XConverter.scala 61:33]
  wire [31:0] fifo_h2c_data_io__in_bits_tuser_mdata; // @[XConverter.scala 61:33]
  wire [5:0] fifo_h2c_data_io__in_bits_tuser_mty; // @[XConverter.scala 61:33]
  wire  fifo_h2c_data_io__in_bits_tuser_zero_byte; // @[XConverter.scala 61:33]
  wire  fifo_h2c_data_io__in_bits_last; // @[XConverter.scala 61:33]
  wire  fifo_h2c_data_io__out_valid; // @[XConverter.scala 61:33]
  wire  fifo_h2c_data_io_in_ready; // @[XConverter.scala 61:33]
  wire  fifo_h2c_data_io_in_valid; // @[XConverter.scala 61:33]
  wire  fifo_h2c_data_io_in_queue_clock; // @[RegSlices.scala 64:35]
  wire  fifo_h2c_data_io_in_queue_reset; // @[RegSlices.scala 64:35]
  wire  fifo_h2c_data_io_in_queue_io_upStream_ready; // @[RegSlices.scala 64:35]
  wire  fifo_h2c_data_io_in_queue_io_upStream_valid; // @[RegSlices.scala 64:35]
  wire [511:0] fifo_h2c_data_io_in_queue_io_upStream_bits_data; // @[RegSlices.scala 64:35]
  wire [31:0] fifo_h2c_data_io_in_queue_io_upStream_bits_tcrc; // @[RegSlices.scala 64:35]
  wire [10:0] fifo_h2c_data_io_in_queue_io_upStream_bits_tuser_qid; // @[RegSlices.scala 64:35]
  wire [2:0] fifo_h2c_data_io_in_queue_io_upStream_bits_tuser_port_id; // @[RegSlices.scala 64:35]
  wire  fifo_h2c_data_io_in_queue_io_upStream_bits_tuser_err; // @[RegSlices.scala 64:35]
  wire [31:0] fifo_h2c_data_io_in_queue_io_upStream_bits_tuser_mdata; // @[RegSlices.scala 64:35]
  wire [5:0] fifo_h2c_data_io_in_queue_io_upStream_bits_tuser_mty; // @[RegSlices.scala 64:35]
  wire  fifo_h2c_data_io_in_queue_io_upStream_bits_tuser_zero_byte; // @[RegSlices.scala 64:35]
  wire  fifo_h2c_data_io_in_queue_io_upStream_bits_last; // @[RegSlices.scala 64:35]
  wire  fifo_h2c_data_io_in_queue_io_downStream_ready; // @[RegSlices.scala 64:35]
  wire  fifo_h2c_data_io_in_queue_io_downStream_valid; // @[RegSlices.scala 64:35]
  wire [511:0] fifo_h2c_data_io_in_queue_io_downStream_bits_data; // @[RegSlices.scala 64:35]
  wire [31:0] fifo_h2c_data_io_in_queue_io_downStream_bits_tcrc; // @[RegSlices.scala 64:35]
  wire [10:0] fifo_h2c_data_io_in_queue_io_downStream_bits_tuser_qid; // @[RegSlices.scala 64:35]
  wire [2:0] fifo_h2c_data_io_in_queue_io_downStream_bits_tuser_port_id; // @[RegSlices.scala 64:35]
  wire  fifo_h2c_data_io_in_queue_io_downStream_bits_tuser_err; // @[RegSlices.scala 64:35]
  wire [31:0] fifo_h2c_data_io_in_queue_io_downStream_bits_tuser_mdata; // @[RegSlices.scala 64:35]
  wire [5:0] fifo_h2c_data_io_in_queue_io_downStream_bits_tuser_mty; // @[RegSlices.scala 64:35]
  wire  fifo_h2c_data_io_in_queue_io_downStream_bits_tuser_zero_byte; // @[RegSlices.scala 64:35]
  wire  fifo_h2c_data_io_in_queue_io_downStream_bits_last; // @[RegSlices.scala 64:35]
  wire  fifo_c2h_data_io__in_clk; // @[XConverter.scala 61:33]
  wire  fifo_c2h_data_io__out_clk; // @[XConverter.scala 61:33]
  wire  fifo_c2h_data_io__rstn; // @[XConverter.scala 61:33]
  wire  fifo_c2h_data_io__in_ready; // @[XConverter.scala 61:33]
  wire  fifo_c2h_data_io__in_valid; // @[XConverter.scala 61:33]
  wire [511:0] fifo_c2h_data_io__in_bits_data; // @[XConverter.scala 61:33]
  wire [31:0] fifo_c2h_data_io__in_bits_tcrc; // @[XConverter.scala 61:33]
  wire  fifo_c2h_data_io__in_bits_ctrl_marker; // @[XConverter.scala 61:33]
  wire [6:0] fifo_c2h_data_io__in_bits_ctrl_ecc; // @[XConverter.scala 61:33]
  wire [31:0] fifo_c2h_data_io__in_bits_ctrl_len; // @[XConverter.scala 61:33]
  wire [2:0] fifo_c2h_data_io__in_bits_ctrl_port_id; // @[XConverter.scala 61:33]
  wire [10:0] fifo_c2h_data_io__in_bits_ctrl_qid; // @[XConverter.scala 61:33]
  wire  fifo_c2h_data_io__in_bits_ctrl_has_cmpt; // @[XConverter.scala 61:33]
  wire  fifo_c2h_data_io__in_bits_last; // @[XConverter.scala 61:33]
  wire [5:0] fifo_c2h_data_io__in_bits_mty; // @[XConverter.scala 61:33]
  wire  fifo_c2h_data_io__out_ready; // @[XConverter.scala 61:33]
  wire  fifo_c2h_data_io__out_valid; // @[XConverter.scala 61:33]
  wire [511:0] fifo_c2h_data_io__out_bits_data; // @[XConverter.scala 61:33]
  wire [31:0] fifo_c2h_data_io__out_bits_tcrc; // @[XConverter.scala 61:33]
  wire  fifo_c2h_data_io__out_bits_ctrl_marker; // @[XConverter.scala 61:33]
  wire [6:0] fifo_c2h_data_io__out_bits_ctrl_ecc; // @[XConverter.scala 61:33]
  wire [31:0] fifo_c2h_data_io__out_bits_ctrl_len; // @[XConverter.scala 61:33]
  wire [2:0] fifo_c2h_data_io__out_bits_ctrl_port_id; // @[XConverter.scala 61:33]
  wire [10:0] fifo_c2h_data_io__out_bits_ctrl_qid; // @[XConverter.scala 61:33]
  wire  fifo_c2h_data_io__out_bits_ctrl_has_cmpt; // @[XConverter.scala 61:33]
  wire  fifo_c2h_data_io__out_bits_last; // @[XConverter.scala 61:33]
  wire [5:0] fifo_c2h_data_io__out_bits_mty; // @[XConverter.scala 61:33]
  wire  fifo_c2h_data_io_out_ready; // @[XConverter.scala 61:33]
  wire  fifo_c2h_data_io_out_valid_0; // @[XConverter.scala 61:33]
  wire  fifo_c2h_data_out_queue_clock; // @[RegSlices.scala 64:35]
  wire  fifo_c2h_data_out_queue_reset; // @[RegSlices.scala 64:35]
  wire  fifo_c2h_data_out_queue_io_upStream_ready; // @[RegSlices.scala 64:35]
  wire  fifo_c2h_data_out_queue_io_upStream_valid; // @[RegSlices.scala 64:35]
  wire [511:0] fifo_c2h_data_out_queue_io_upStream_bits_data; // @[RegSlices.scala 64:35]
  wire [31:0] fifo_c2h_data_out_queue_io_upStream_bits_tcrc; // @[RegSlices.scala 64:35]
  wire  fifo_c2h_data_out_queue_io_upStream_bits_ctrl_marker; // @[RegSlices.scala 64:35]
  wire [6:0] fifo_c2h_data_out_queue_io_upStream_bits_ctrl_ecc; // @[RegSlices.scala 64:35]
  wire [31:0] fifo_c2h_data_out_queue_io_upStream_bits_ctrl_len; // @[RegSlices.scala 64:35]
  wire [2:0] fifo_c2h_data_out_queue_io_upStream_bits_ctrl_port_id; // @[RegSlices.scala 64:35]
  wire [10:0] fifo_c2h_data_out_queue_io_upStream_bits_ctrl_qid; // @[RegSlices.scala 64:35]
  wire  fifo_c2h_data_out_queue_io_upStream_bits_ctrl_has_cmpt; // @[RegSlices.scala 64:35]
  wire  fifo_c2h_data_out_queue_io_upStream_bits_last; // @[RegSlices.scala 64:35]
  wire [5:0] fifo_c2h_data_out_queue_io_upStream_bits_mty; // @[RegSlices.scala 64:35]
  wire  fifo_c2h_data_out_queue_io_downStream_ready; // @[RegSlices.scala 64:35]
  wire  fifo_c2h_data_out_queue_io_downStream_valid; // @[RegSlices.scala 64:35]
  wire [511:0] fifo_c2h_data_out_queue_io_downStream_bits_data; // @[RegSlices.scala 64:35]
  wire [31:0] fifo_c2h_data_out_queue_io_downStream_bits_tcrc; // @[RegSlices.scala 64:35]
  wire  fifo_c2h_data_out_queue_io_downStream_bits_ctrl_marker; // @[RegSlices.scala 64:35]
  wire [6:0] fifo_c2h_data_out_queue_io_downStream_bits_ctrl_ecc; // @[RegSlices.scala 64:35]
  wire [31:0] fifo_c2h_data_out_queue_io_downStream_bits_ctrl_len; // @[RegSlices.scala 64:35]
  wire [2:0] fifo_c2h_data_out_queue_io_downStream_bits_ctrl_port_id; // @[RegSlices.scala 64:35]
  wire [10:0] fifo_c2h_data_out_queue_io_downStream_bits_ctrl_qid; // @[RegSlices.scala 64:35]
  wire  fifo_c2h_data_out_queue_io_downStream_bits_ctrl_has_cmpt; // @[RegSlices.scala 64:35]
  wire  fifo_c2h_data_out_queue_io_downStream_bits_last; // @[RegSlices.scala 64:35]
  wire [5:0] fifo_c2h_data_out_queue_io_downStream_bits_mty; // @[RegSlices.scala 64:35]
  wire  fifo_h2c_cmd_io__in_clk; // @[XConverter.scala 61:33]
  wire  fifo_h2c_cmd_io__out_clk; // @[XConverter.scala 61:33]
  wire  fifo_h2c_cmd_io__rstn; // @[XConverter.scala 61:33]
  wire  fifo_h2c_cmd_io__in_ready; // @[XConverter.scala 61:33]
  wire  fifo_h2c_cmd_io__in_valid; // @[XConverter.scala 61:33]
  wire [63:0] fifo_h2c_cmd_io__in_bits_addr; // @[XConverter.scala 61:33]
  wire [31:0] fifo_h2c_cmd_io__in_bits_len; // @[XConverter.scala 61:33]
  wire  fifo_h2c_cmd_io__in_bits_eop; // @[XConverter.scala 61:33]
  wire  fifo_h2c_cmd_io__in_bits_sop; // @[XConverter.scala 61:33]
  wire  fifo_h2c_cmd_io__in_bits_mrkr_req; // @[XConverter.scala 61:33]
  wire  fifo_h2c_cmd_io__in_bits_sdi; // @[XConverter.scala 61:33]
  wire [10:0] fifo_h2c_cmd_io__in_bits_qid; // @[XConverter.scala 61:33]
  wire  fifo_h2c_cmd_io__in_bits_error; // @[XConverter.scala 61:33]
  wire [7:0] fifo_h2c_cmd_io__in_bits_func; // @[XConverter.scala 61:33]
  wire [15:0] fifo_h2c_cmd_io__in_bits_cidx; // @[XConverter.scala 61:33]
  wire [2:0] fifo_h2c_cmd_io__in_bits_port_id; // @[XConverter.scala 61:33]
  wire  fifo_h2c_cmd_io__in_bits_no_dma; // @[XConverter.scala 61:33]
  wire  fifo_h2c_cmd_io__out_ready; // @[XConverter.scala 61:33]
  wire  fifo_h2c_cmd_io__out_valid; // @[XConverter.scala 61:33]
  wire [63:0] fifo_h2c_cmd_io__out_bits_addr; // @[XConverter.scala 61:33]
  wire [31:0] fifo_h2c_cmd_io__out_bits_len; // @[XConverter.scala 61:33]
  wire  fifo_h2c_cmd_io__out_bits_eop; // @[XConverter.scala 61:33]
  wire  fifo_h2c_cmd_io__out_bits_sop; // @[XConverter.scala 61:33]
  wire  fifo_h2c_cmd_io__out_bits_mrkr_req; // @[XConverter.scala 61:33]
  wire  fifo_h2c_cmd_io__out_bits_sdi; // @[XConverter.scala 61:33]
  wire [10:0] fifo_h2c_cmd_io__out_bits_qid; // @[XConverter.scala 61:33]
  wire  fifo_h2c_cmd_io__out_bits_error; // @[XConverter.scala 61:33]
  wire [7:0] fifo_h2c_cmd_io__out_bits_func; // @[XConverter.scala 61:33]
  wire [15:0] fifo_h2c_cmd_io__out_bits_cidx; // @[XConverter.scala 61:33]
  wire [2:0] fifo_h2c_cmd_io__out_bits_port_id; // @[XConverter.scala 61:33]
  wire  fifo_h2c_cmd_io__out_bits_no_dma; // @[XConverter.scala 61:33]
  wire  fifo_h2c_cmd_io_out_valid; // @[XConverter.scala 61:33]
  wire  fifo_h2c_cmd_io_out_ready_1; // @[XConverter.scala 61:33]
  wire  fifo_h2c_cmd_out_queue_clock; // @[RegSlices.scala 64:35]
  wire  fifo_h2c_cmd_out_queue_reset; // @[RegSlices.scala 64:35]
  wire  fifo_h2c_cmd_out_queue_io_upStream_ready; // @[RegSlices.scala 64:35]
  wire  fifo_h2c_cmd_out_queue_io_upStream_valid; // @[RegSlices.scala 64:35]
  wire [63:0] fifo_h2c_cmd_out_queue_io_upStream_bits_addr; // @[RegSlices.scala 64:35]
  wire [31:0] fifo_h2c_cmd_out_queue_io_upStream_bits_len; // @[RegSlices.scala 64:35]
  wire  fifo_h2c_cmd_out_queue_io_upStream_bits_eop; // @[RegSlices.scala 64:35]
  wire  fifo_h2c_cmd_out_queue_io_upStream_bits_sop; // @[RegSlices.scala 64:35]
  wire  fifo_h2c_cmd_out_queue_io_upStream_bits_mrkr_req; // @[RegSlices.scala 64:35]
  wire  fifo_h2c_cmd_out_queue_io_upStream_bits_sdi; // @[RegSlices.scala 64:35]
  wire [10:0] fifo_h2c_cmd_out_queue_io_upStream_bits_qid; // @[RegSlices.scala 64:35]
  wire  fifo_h2c_cmd_out_queue_io_upStream_bits_error; // @[RegSlices.scala 64:35]
  wire [7:0] fifo_h2c_cmd_out_queue_io_upStream_bits_func; // @[RegSlices.scala 64:35]
  wire [15:0] fifo_h2c_cmd_out_queue_io_upStream_bits_cidx; // @[RegSlices.scala 64:35]
  wire [2:0] fifo_h2c_cmd_out_queue_io_upStream_bits_port_id; // @[RegSlices.scala 64:35]
  wire  fifo_h2c_cmd_out_queue_io_upStream_bits_no_dma; // @[RegSlices.scala 64:35]
  wire  fifo_h2c_cmd_out_queue_io_downStream_ready; // @[RegSlices.scala 64:35]
  wire  fifo_h2c_cmd_out_queue_io_downStream_valid; // @[RegSlices.scala 64:35]
  wire [63:0] fifo_h2c_cmd_out_queue_io_downStream_bits_addr; // @[RegSlices.scala 64:35]
  wire [31:0] fifo_h2c_cmd_out_queue_io_downStream_bits_len; // @[RegSlices.scala 64:35]
  wire  fifo_h2c_cmd_out_queue_io_downStream_bits_eop; // @[RegSlices.scala 64:35]
  wire  fifo_h2c_cmd_out_queue_io_downStream_bits_sop; // @[RegSlices.scala 64:35]
  wire  fifo_h2c_cmd_out_queue_io_downStream_bits_mrkr_req; // @[RegSlices.scala 64:35]
  wire  fifo_h2c_cmd_out_queue_io_downStream_bits_sdi; // @[RegSlices.scala 64:35]
  wire [10:0] fifo_h2c_cmd_out_queue_io_downStream_bits_qid; // @[RegSlices.scala 64:35]
  wire  fifo_h2c_cmd_out_queue_io_downStream_bits_error; // @[RegSlices.scala 64:35]
  wire [7:0] fifo_h2c_cmd_out_queue_io_downStream_bits_func; // @[RegSlices.scala 64:35]
  wire [15:0] fifo_h2c_cmd_out_queue_io_downStream_bits_cidx; // @[RegSlices.scala 64:35]
  wire [2:0] fifo_h2c_cmd_out_queue_io_downStream_bits_port_id; // @[RegSlices.scala 64:35]
  wire  fifo_h2c_cmd_out_queue_io_downStream_bits_no_dma; // @[RegSlices.scala 64:35]
  wire  fifo_c2h_cmd_io_in_clk; // @[XConverter.scala 61:33]
  wire  fifo_c2h_cmd_io_out_clk; // @[XConverter.scala 61:33]
  wire  fifo_c2h_cmd_io_rstn; // @[XConverter.scala 61:33]
  wire  fifo_c2h_cmd_io_in_ready; // @[XConverter.scala 61:33]
  wire  fifo_c2h_cmd_io_in_valid; // @[XConverter.scala 61:33]
  wire [63:0] fifo_c2h_cmd_io_in_bits_addr; // @[XConverter.scala 61:33]
  wire [10:0] fifo_c2h_cmd_io_in_bits_qid; // @[XConverter.scala 61:33]
  wire  fifo_c2h_cmd_io_in_bits_error; // @[XConverter.scala 61:33]
  wire [7:0] fifo_c2h_cmd_io_in_bits_func; // @[XConverter.scala 61:33]
  wire [2:0] fifo_c2h_cmd_io_in_bits_port_id; // @[XConverter.scala 61:33]
  wire [6:0] fifo_c2h_cmd_io_in_bits_pfch_tag; // @[XConverter.scala 61:33]
  wire [31:0] fifo_c2h_cmd_io_in_bits_len; // @[XConverter.scala 61:33]
  wire  fifo_c2h_cmd_io_out_ready; // @[XConverter.scala 61:33]
  wire  fifo_c2h_cmd_io_out_valid; // @[XConverter.scala 61:33]
  wire [63:0] fifo_c2h_cmd_io_out_bits_addr; // @[XConverter.scala 61:33]
  wire [10:0] fifo_c2h_cmd_io_out_bits_qid; // @[XConverter.scala 61:33]
  wire  fifo_c2h_cmd_io_out_bits_error; // @[XConverter.scala 61:33]
  wire [7:0] fifo_c2h_cmd_io_out_bits_func; // @[XConverter.scala 61:33]
  wire [2:0] fifo_c2h_cmd_io_out_bits_port_id; // @[XConverter.scala 61:33]
  wire [6:0] fifo_c2h_cmd_io_out_bits_pfch_tag; // @[XConverter.scala 61:33]
  wire [31:0] fifo_c2h_cmd_io_out_bits_len; // @[XConverter.scala 61:33]
  wire  fifo_c2h_cmd_io_out_ready_0; // @[XConverter.scala 61:33]
  wire  fifo_c2h_cmd_io_out_valid_1; // @[XConverter.scala 61:33]
  wire  fifo_c2h_cmd_out_queue_clock; // @[RegSlices.scala 64:35]
  wire  fifo_c2h_cmd_out_queue_reset; // @[RegSlices.scala 64:35]
  wire  fifo_c2h_cmd_out_queue_io_upStream_ready; // @[RegSlices.scala 64:35]
  wire  fifo_c2h_cmd_out_queue_io_upStream_valid; // @[RegSlices.scala 64:35]
  wire [63:0] fifo_c2h_cmd_out_queue_io_upStream_bits_addr; // @[RegSlices.scala 64:35]
  wire [10:0] fifo_c2h_cmd_out_queue_io_upStream_bits_qid; // @[RegSlices.scala 64:35]
  wire  fifo_c2h_cmd_out_queue_io_upStream_bits_error; // @[RegSlices.scala 64:35]
  wire [7:0] fifo_c2h_cmd_out_queue_io_upStream_bits_func; // @[RegSlices.scala 64:35]
  wire [2:0] fifo_c2h_cmd_out_queue_io_upStream_bits_port_id; // @[RegSlices.scala 64:35]
  wire [6:0] fifo_c2h_cmd_out_queue_io_upStream_bits_pfch_tag; // @[RegSlices.scala 64:35]
  wire [31:0] fifo_c2h_cmd_out_queue_io_upStream_bits_len; // @[RegSlices.scala 64:35]
  wire  fifo_c2h_cmd_out_queue_io_downStream_ready; // @[RegSlices.scala 64:35]
  wire  fifo_c2h_cmd_out_queue_io_downStream_valid; // @[RegSlices.scala 64:35]
  wire [63:0] fifo_c2h_cmd_out_queue_io_downStream_bits_addr; // @[RegSlices.scala 64:35]
  wire [10:0] fifo_c2h_cmd_out_queue_io_downStream_bits_qid; // @[RegSlices.scala 64:35]
  wire  fifo_c2h_cmd_out_queue_io_downStream_bits_error; // @[RegSlices.scala 64:35]
  wire [7:0] fifo_c2h_cmd_out_queue_io_downStream_bits_func; // @[RegSlices.scala 64:35]
  wire [2:0] fifo_c2h_cmd_out_queue_io_downStream_bits_port_id; // @[RegSlices.scala 64:35]
  wire [6:0] fifo_c2h_cmd_out_queue_io_downStream_bits_pfch_tag; // @[RegSlices.scala 64:35]
  wire [31:0] fifo_c2h_cmd_out_queue_io_downStream_bits_len; // @[RegSlices.scala 64:35]
  wire  check_c2h_clock; // @[QDMADynamic.scala 62:95]
  wire  check_c2h_reset; // @[QDMADynamic.scala 62:95]
  wire  check_c2h_io_in_ready; // @[QDMADynamic.scala 62:95]
  wire  check_c2h_io_in_valid; // @[QDMADynamic.scala 62:95]
  wire [63:0] check_c2h_io_in_bits_addr; // @[QDMADynamic.scala 62:95]
  wire [10:0] check_c2h_io_in_bits_qid; // @[QDMADynamic.scala 62:95]
  wire  check_c2h_io_in_bits_error; // @[QDMADynamic.scala 62:95]
  wire [7:0] check_c2h_io_in_bits_func; // @[QDMADynamic.scala 62:95]
  wire [2:0] check_c2h_io_in_bits_port_id; // @[QDMADynamic.scala 62:95]
  wire [6:0] check_c2h_io_in_bits_pfch_tag; // @[QDMADynamic.scala 62:95]
  wire [31:0] check_c2h_io_in_bits_len; // @[QDMADynamic.scala 62:95]
  wire  check_c2h_io_out_ready; // @[QDMADynamic.scala 62:95]
  wire  check_c2h_io_out_valid; // @[QDMADynamic.scala 62:95]
  wire [63:0] check_c2h_io_out_bits_addr; // @[QDMADynamic.scala 62:95]
  wire [10:0] check_c2h_io_out_bits_qid; // @[QDMADynamic.scala 62:95]
  wire  check_c2h_io_out_bits_error; // @[QDMADynamic.scala 62:95]
  wire [7:0] check_c2h_io_out_bits_func; // @[QDMADynamic.scala 62:95]
  wire [2:0] check_c2h_io_out_bits_port_id; // @[QDMADynamic.scala 62:95]
  wire [6:0] check_c2h_io_out_bits_pfch_tag; // @[QDMADynamic.scala 62:95]
  wire [31:0] check_c2h_io_out_bits_len; // @[QDMADynamic.scala 62:95]
  wire  check_c2h_io_in_queue_clock; // @[RegSlices.scala 64:35]
  wire  check_c2h_io_in_queue_reset; // @[RegSlices.scala 64:35]
  wire  check_c2h_io_in_queue_io_upStream_ready; // @[RegSlices.scala 64:35]
  wire  check_c2h_io_in_queue_io_upStream_valid; // @[RegSlices.scala 64:35]
  wire [63:0] check_c2h_io_in_queue_io_upStream_bits_addr; // @[RegSlices.scala 64:35]
  wire [10:0] check_c2h_io_in_queue_io_upStream_bits_qid; // @[RegSlices.scala 64:35]
  wire  check_c2h_io_in_queue_io_upStream_bits_error; // @[RegSlices.scala 64:35]
  wire [7:0] check_c2h_io_in_queue_io_upStream_bits_func; // @[RegSlices.scala 64:35]
  wire [2:0] check_c2h_io_in_queue_io_upStream_bits_port_id; // @[RegSlices.scala 64:35]
  wire [6:0] check_c2h_io_in_queue_io_upStream_bits_pfch_tag; // @[RegSlices.scala 64:35]
  wire [31:0] check_c2h_io_in_queue_io_upStream_bits_len; // @[RegSlices.scala 64:35]
  wire  check_c2h_io_in_queue_io_downStream_ready; // @[RegSlices.scala 64:35]
  wire  check_c2h_io_in_queue_io_downStream_valid; // @[RegSlices.scala 64:35]
  wire [63:0] check_c2h_io_in_queue_io_downStream_bits_addr; // @[RegSlices.scala 64:35]
  wire [10:0] check_c2h_io_in_queue_io_downStream_bits_qid; // @[RegSlices.scala 64:35]
  wire  check_c2h_io_in_queue_io_downStream_bits_error; // @[RegSlices.scala 64:35]
  wire [7:0] check_c2h_io_in_queue_io_downStream_bits_func; // @[RegSlices.scala 64:35]
  wire [2:0] check_c2h_io_in_queue_io_downStream_bits_port_id; // @[RegSlices.scala 64:35]
  wire [6:0] check_c2h_io_in_queue_io_downStream_bits_pfch_tag; // @[RegSlices.scala 64:35]
  wire [31:0] check_c2h_io_in_queue_io_downStream_bits_len; // @[RegSlices.scala 64:35]
  wire  check_h2c_clock; // @[QDMADynamic.scala 64:95]
  wire  check_h2c_reset; // @[QDMADynamic.scala 64:95]
  wire  check_h2c_io_in_ready; // @[QDMADynamic.scala 64:95]
  wire  check_h2c_io_in_valid; // @[QDMADynamic.scala 64:95]
  wire [63:0] check_h2c_io_in_bits_addr; // @[QDMADynamic.scala 64:95]
  wire [31:0] check_h2c_io_in_bits_len; // @[QDMADynamic.scala 64:95]
  wire  check_h2c_io_in_bits_eop; // @[QDMADynamic.scala 64:95]
  wire  check_h2c_io_in_bits_sop; // @[QDMADynamic.scala 64:95]
  wire  check_h2c_io_in_bits_mrkr_req; // @[QDMADynamic.scala 64:95]
  wire  check_h2c_io_in_bits_sdi; // @[QDMADynamic.scala 64:95]
  wire [10:0] check_h2c_io_in_bits_qid; // @[QDMADynamic.scala 64:95]
  wire  check_h2c_io_in_bits_error; // @[QDMADynamic.scala 64:95]
  wire [7:0] check_h2c_io_in_bits_func; // @[QDMADynamic.scala 64:95]
  wire [15:0] check_h2c_io_in_bits_cidx; // @[QDMADynamic.scala 64:95]
  wire [2:0] check_h2c_io_in_bits_port_id; // @[QDMADynamic.scala 64:95]
  wire  check_h2c_io_in_bits_no_dma; // @[QDMADynamic.scala 64:95]
  wire  check_h2c_io_out_ready; // @[QDMADynamic.scala 64:95]
  wire  check_h2c_io_out_valid; // @[QDMADynamic.scala 64:95]
  wire [63:0] check_h2c_io_out_bits_addr; // @[QDMADynamic.scala 64:95]
  wire [31:0] check_h2c_io_out_bits_len; // @[QDMADynamic.scala 64:95]
  wire  check_h2c_io_out_bits_eop; // @[QDMADynamic.scala 64:95]
  wire  check_h2c_io_out_bits_sop; // @[QDMADynamic.scala 64:95]
  wire  check_h2c_io_out_bits_mrkr_req; // @[QDMADynamic.scala 64:95]
  wire  check_h2c_io_out_bits_sdi; // @[QDMADynamic.scala 64:95]
  wire [10:0] check_h2c_io_out_bits_qid; // @[QDMADynamic.scala 64:95]
  wire  check_h2c_io_out_bits_error; // @[QDMADynamic.scala 64:95]
  wire [7:0] check_h2c_io_out_bits_func; // @[QDMADynamic.scala 64:95]
  wire [15:0] check_h2c_io_out_bits_cidx; // @[QDMADynamic.scala 64:95]
  wire [2:0] check_h2c_io_out_bits_port_id; // @[QDMADynamic.scala 64:95]
  wire  check_h2c_io_out_bits_no_dma; // @[QDMADynamic.scala 64:95]
  wire  check_h2c_io_in_queue_clock; // @[RegSlices.scala 64:35]
  wire  check_h2c_io_in_queue_reset; // @[RegSlices.scala 64:35]
  wire  check_h2c_io_in_queue_io_upStream_ready; // @[RegSlices.scala 64:35]
  wire  check_h2c_io_in_queue_io_upStream_valid; // @[RegSlices.scala 64:35]
  wire [63:0] check_h2c_io_in_queue_io_upStream_bits_addr; // @[RegSlices.scala 64:35]
  wire [31:0] check_h2c_io_in_queue_io_upStream_bits_len; // @[RegSlices.scala 64:35]
  wire  check_h2c_io_in_queue_io_upStream_bits_eop; // @[RegSlices.scala 64:35]
  wire  check_h2c_io_in_queue_io_upStream_bits_sop; // @[RegSlices.scala 64:35]
  wire  check_h2c_io_in_queue_io_upStream_bits_mrkr_req; // @[RegSlices.scala 64:35]
  wire  check_h2c_io_in_queue_io_upStream_bits_sdi; // @[RegSlices.scala 64:35]
  wire [10:0] check_h2c_io_in_queue_io_upStream_bits_qid; // @[RegSlices.scala 64:35]
  wire  check_h2c_io_in_queue_io_upStream_bits_error; // @[RegSlices.scala 64:35]
  wire [7:0] check_h2c_io_in_queue_io_upStream_bits_func; // @[RegSlices.scala 64:35]
  wire [15:0] check_h2c_io_in_queue_io_upStream_bits_cidx; // @[RegSlices.scala 64:35]
  wire [2:0] check_h2c_io_in_queue_io_upStream_bits_port_id; // @[RegSlices.scala 64:35]
  wire  check_h2c_io_in_queue_io_upStream_bits_no_dma; // @[RegSlices.scala 64:35]
  wire  check_h2c_io_in_queue_io_downStream_ready; // @[RegSlices.scala 64:35]
  wire  check_h2c_io_in_queue_io_downStream_valid; // @[RegSlices.scala 64:35]
  wire [63:0] check_h2c_io_in_queue_io_downStream_bits_addr; // @[RegSlices.scala 64:35]
  wire [31:0] check_h2c_io_in_queue_io_downStream_bits_len; // @[RegSlices.scala 64:35]
  wire  check_h2c_io_in_queue_io_downStream_bits_eop; // @[RegSlices.scala 64:35]
  wire  check_h2c_io_in_queue_io_downStream_bits_sop; // @[RegSlices.scala 64:35]
  wire  check_h2c_io_in_queue_io_downStream_bits_mrkr_req; // @[RegSlices.scala 64:35]
  wire  check_h2c_io_in_queue_io_downStream_bits_sdi; // @[RegSlices.scala 64:35]
  wire [10:0] check_h2c_io_in_queue_io_downStream_bits_qid; // @[RegSlices.scala 64:35]
  wire  check_h2c_io_in_queue_io_downStream_bits_error; // @[RegSlices.scala 64:35]
  wire [7:0] check_h2c_io_in_queue_io_downStream_bits_func; // @[RegSlices.scala 64:35]
  wire [15:0] check_h2c_io_in_queue_io_downStream_bits_cidx; // @[RegSlices.scala 64:35]
  wire [2:0] check_h2c_io_in_queue_io_downStream_bits_port_id; // @[RegSlices.scala 64:35]
  wire  check_h2c_io_in_queue_io_downStream_bits_no_dma; // @[RegSlices.scala 64:35]
  wire  tlb_clock; // @[QDMADynamic.scala 67:71]
  wire  tlb_reset; // @[QDMADynamic.scala 67:71]
  wire  tlb_io__wr_tlb_ready; // @[QDMADynamic.scala 67:71]
  wire  tlb_io__wr_tlb_valid; // @[QDMADynamic.scala 67:71]
  wire [31:0] tlb_io__wr_tlb_bits_vaddr_high; // @[QDMADynamic.scala 67:71]
  wire [31:0] tlb_io__wr_tlb_bits_vaddr_low; // @[QDMADynamic.scala 67:71]
  wire [31:0] tlb_io__wr_tlb_bits_paddr_high; // @[QDMADynamic.scala 67:71]
  wire [31:0] tlb_io__wr_tlb_bits_paddr_low; // @[QDMADynamic.scala 67:71]
  wire  tlb_io__wr_tlb_bits_is_base; // @[QDMADynamic.scala 67:71]
  wire  tlb_io__h2c_in_ready; // @[QDMADynamic.scala 67:71]
  wire  tlb_io__h2c_in_valid; // @[QDMADynamic.scala 67:71]
  wire [63:0] tlb_io__h2c_in_bits_addr; // @[QDMADynamic.scala 67:71]
  wire [31:0] tlb_io__h2c_in_bits_len; // @[QDMADynamic.scala 67:71]
  wire  tlb_io__h2c_in_bits_eop; // @[QDMADynamic.scala 67:71]
  wire  tlb_io__h2c_in_bits_sop; // @[QDMADynamic.scala 67:71]
  wire  tlb_io__h2c_in_bits_mrkr_req; // @[QDMADynamic.scala 67:71]
  wire  tlb_io__h2c_in_bits_sdi; // @[QDMADynamic.scala 67:71]
  wire [10:0] tlb_io__h2c_in_bits_qid; // @[QDMADynamic.scala 67:71]
  wire  tlb_io__h2c_in_bits_error; // @[QDMADynamic.scala 67:71]
  wire [7:0] tlb_io__h2c_in_bits_func; // @[QDMADynamic.scala 67:71]
  wire [15:0] tlb_io__h2c_in_bits_cidx; // @[QDMADynamic.scala 67:71]
  wire [2:0] tlb_io__h2c_in_bits_port_id; // @[QDMADynamic.scala 67:71]
  wire  tlb_io__h2c_in_bits_no_dma; // @[QDMADynamic.scala 67:71]
  wire  tlb_io__c2h_in_ready; // @[QDMADynamic.scala 67:71]
  wire  tlb_io__c2h_in_valid; // @[QDMADynamic.scala 67:71]
  wire [63:0] tlb_io__c2h_in_bits_addr; // @[QDMADynamic.scala 67:71]
  wire [10:0] tlb_io__c2h_in_bits_qid; // @[QDMADynamic.scala 67:71]
  wire  tlb_io__c2h_in_bits_error; // @[QDMADynamic.scala 67:71]
  wire [7:0] tlb_io__c2h_in_bits_func; // @[QDMADynamic.scala 67:71]
  wire [2:0] tlb_io__c2h_in_bits_port_id; // @[QDMADynamic.scala 67:71]
  wire [6:0] tlb_io__c2h_in_bits_pfch_tag; // @[QDMADynamic.scala 67:71]
  wire [31:0] tlb_io__c2h_in_bits_len; // @[QDMADynamic.scala 67:71]
  wire  tlb_io__h2c_out_ready; // @[QDMADynamic.scala 67:71]
  wire  tlb_io__h2c_out_valid; // @[QDMADynamic.scala 67:71]
  wire [63:0] tlb_io__h2c_out_bits_addr; // @[QDMADynamic.scala 67:71]
  wire [31:0] tlb_io__h2c_out_bits_len; // @[QDMADynamic.scala 67:71]
  wire  tlb_io__h2c_out_bits_eop; // @[QDMADynamic.scala 67:71]
  wire  tlb_io__h2c_out_bits_sop; // @[QDMADynamic.scala 67:71]
  wire  tlb_io__h2c_out_bits_mrkr_req; // @[QDMADynamic.scala 67:71]
  wire  tlb_io__h2c_out_bits_sdi; // @[QDMADynamic.scala 67:71]
  wire [10:0] tlb_io__h2c_out_bits_qid; // @[QDMADynamic.scala 67:71]
  wire  tlb_io__h2c_out_bits_error; // @[QDMADynamic.scala 67:71]
  wire [7:0] tlb_io__h2c_out_bits_func; // @[QDMADynamic.scala 67:71]
  wire [15:0] tlb_io__h2c_out_bits_cidx; // @[QDMADynamic.scala 67:71]
  wire [2:0] tlb_io__h2c_out_bits_port_id; // @[QDMADynamic.scala 67:71]
  wire  tlb_io__h2c_out_bits_no_dma; // @[QDMADynamic.scala 67:71]
  wire  tlb_io__c2h_out_ready; // @[QDMADynamic.scala 67:71]
  wire  tlb_io__c2h_out_valid; // @[QDMADynamic.scala 67:71]
  wire [63:0] tlb_io__c2h_out_bits_addr; // @[QDMADynamic.scala 67:71]
  wire [10:0] tlb_io__c2h_out_bits_qid; // @[QDMADynamic.scala 67:71]
  wire  tlb_io__c2h_out_bits_error; // @[QDMADynamic.scala 67:71]
  wire [7:0] tlb_io__c2h_out_bits_func; // @[QDMADynamic.scala 67:71]
  wire [2:0] tlb_io__c2h_out_bits_port_id; // @[QDMADynamic.scala 67:71]
  wire [6:0] tlb_io__c2h_out_bits_pfch_tag; // @[QDMADynamic.scala 67:71]
  wire [31:0] tlb_io__c2h_out_bits_len; // @[QDMADynamic.scala 67:71]
  wire [31:0] tlb_io__tlb_miss_count; // @[QDMADynamic.scala 67:71]
  wire [31:0] tlb_io_tlb_miss_count; // @[QDMADynamic.scala 67:71]
  wire  tlb_io_h2c_in_queue_clock; // @[RegSlices.scala 64:35]
  wire  tlb_io_h2c_in_queue_reset; // @[RegSlices.scala 64:35]
  wire  tlb_io_h2c_in_queue_io_upStream_ready; // @[RegSlices.scala 64:35]
  wire  tlb_io_h2c_in_queue_io_upStream_valid; // @[RegSlices.scala 64:35]
  wire [63:0] tlb_io_h2c_in_queue_io_upStream_bits_addr; // @[RegSlices.scala 64:35]
  wire [31:0] tlb_io_h2c_in_queue_io_upStream_bits_len; // @[RegSlices.scala 64:35]
  wire  tlb_io_h2c_in_queue_io_upStream_bits_eop; // @[RegSlices.scala 64:35]
  wire  tlb_io_h2c_in_queue_io_upStream_bits_sop; // @[RegSlices.scala 64:35]
  wire  tlb_io_h2c_in_queue_io_upStream_bits_mrkr_req; // @[RegSlices.scala 64:35]
  wire  tlb_io_h2c_in_queue_io_upStream_bits_sdi; // @[RegSlices.scala 64:35]
  wire [10:0] tlb_io_h2c_in_queue_io_upStream_bits_qid; // @[RegSlices.scala 64:35]
  wire  tlb_io_h2c_in_queue_io_upStream_bits_error; // @[RegSlices.scala 64:35]
  wire [7:0] tlb_io_h2c_in_queue_io_upStream_bits_func; // @[RegSlices.scala 64:35]
  wire [15:0] tlb_io_h2c_in_queue_io_upStream_bits_cidx; // @[RegSlices.scala 64:35]
  wire [2:0] tlb_io_h2c_in_queue_io_upStream_bits_port_id; // @[RegSlices.scala 64:35]
  wire  tlb_io_h2c_in_queue_io_upStream_bits_no_dma; // @[RegSlices.scala 64:35]
  wire  tlb_io_h2c_in_queue_io_downStream_ready; // @[RegSlices.scala 64:35]
  wire  tlb_io_h2c_in_queue_io_downStream_valid; // @[RegSlices.scala 64:35]
  wire [63:0] tlb_io_h2c_in_queue_io_downStream_bits_addr; // @[RegSlices.scala 64:35]
  wire [31:0] tlb_io_h2c_in_queue_io_downStream_bits_len; // @[RegSlices.scala 64:35]
  wire  tlb_io_h2c_in_queue_io_downStream_bits_eop; // @[RegSlices.scala 64:35]
  wire  tlb_io_h2c_in_queue_io_downStream_bits_sop; // @[RegSlices.scala 64:35]
  wire  tlb_io_h2c_in_queue_io_downStream_bits_mrkr_req; // @[RegSlices.scala 64:35]
  wire  tlb_io_h2c_in_queue_io_downStream_bits_sdi; // @[RegSlices.scala 64:35]
  wire [10:0] tlb_io_h2c_in_queue_io_downStream_bits_qid; // @[RegSlices.scala 64:35]
  wire  tlb_io_h2c_in_queue_io_downStream_bits_error; // @[RegSlices.scala 64:35]
  wire [7:0] tlb_io_h2c_in_queue_io_downStream_bits_func; // @[RegSlices.scala 64:35]
  wire [15:0] tlb_io_h2c_in_queue_io_downStream_bits_cidx; // @[RegSlices.scala 64:35]
  wire [2:0] tlb_io_h2c_in_queue_io_downStream_bits_port_id; // @[RegSlices.scala 64:35]
  wire  tlb_io_h2c_in_queue_io_downStream_bits_no_dma; // @[RegSlices.scala 64:35]
  wire  tlb_io_c2h_in_queue_clock; // @[RegSlices.scala 64:35]
  wire  tlb_io_c2h_in_queue_reset; // @[RegSlices.scala 64:35]
  wire  tlb_io_c2h_in_queue_io_upStream_ready; // @[RegSlices.scala 64:35]
  wire  tlb_io_c2h_in_queue_io_upStream_valid; // @[RegSlices.scala 64:35]
  wire [63:0] tlb_io_c2h_in_queue_io_upStream_bits_addr; // @[RegSlices.scala 64:35]
  wire [10:0] tlb_io_c2h_in_queue_io_upStream_bits_qid; // @[RegSlices.scala 64:35]
  wire  tlb_io_c2h_in_queue_io_upStream_bits_error; // @[RegSlices.scala 64:35]
  wire [7:0] tlb_io_c2h_in_queue_io_upStream_bits_func; // @[RegSlices.scala 64:35]
  wire [2:0] tlb_io_c2h_in_queue_io_upStream_bits_port_id; // @[RegSlices.scala 64:35]
  wire [6:0] tlb_io_c2h_in_queue_io_upStream_bits_pfch_tag; // @[RegSlices.scala 64:35]
  wire [31:0] tlb_io_c2h_in_queue_io_upStream_bits_len; // @[RegSlices.scala 64:35]
  wire  tlb_io_c2h_in_queue_io_downStream_ready; // @[RegSlices.scala 64:35]
  wire  tlb_io_c2h_in_queue_io_downStream_valid; // @[RegSlices.scala 64:35]
  wire [63:0] tlb_io_c2h_in_queue_io_downStream_bits_addr; // @[RegSlices.scala 64:35]
  wire [10:0] tlb_io_c2h_in_queue_io_downStream_bits_qid; // @[RegSlices.scala 64:35]
  wire  tlb_io_c2h_in_queue_io_downStream_bits_error; // @[RegSlices.scala 64:35]
  wire [7:0] tlb_io_c2h_in_queue_io_downStream_bits_func; // @[RegSlices.scala 64:35]
  wire [2:0] tlb_io_c2h_in_queue_io_downStream_bits_port_id; // @[RegSlices.scala 64:35]
  wire [6:0] tlb_io_c2h_in_queue_io_downStream_bits_pfch_tag; // @[RegSlices.scala 64:35]
  wire [31:0] tlb_io_c2h_in_queue_io_downStream_bits_len; // @[RegSlices.scala 64:35]
  wire  fifo_h2c_cmd_io_in_queue_clock; // @[RegSlices.scala 64:35]
  wire  fifo_h2c_cmd_io_in_queue_reset; // @[RegSlices.scala 64:35]
  wire  fifo_h2c_cmd_io_in_queue_io_upStream_ready; // @[RegSlices.scala 64:35]
  wire  fifo_h2c_cmd_io_in_queue_io_upStream_valid; // @[RegSlices.scala 64:35]
  wire [63:0] fifo_h2c_cmd_io_in_queue_io_upStream_bits_addr; // @[RegSlices.scala 64:35]
  wire [31:0] fifo_h2c_cmd_io_in_queue_io_upStream_bits_len; // @[RegSlices.scala 64:35]
  wire  fifo_h2c_cmd_io_in_queue_io_upStream_bits_eop; // @[RegSlices.scala 64:35]
  wire  fifo_h2c_cmd_io_in_queue_io_upStream_bits_sop; // @[RegSlices.scala 64:35]
  wire  fifo_h2c_cmd_io_in_queue_io_upStream_bits_mrkr_req; // @[RegSlices.scala 64:35]
  wire  fifo_h2c_cmd_io_in_queue_io_upStream_bits_sdi; // @[RegSlices.scala 64:35]
  wire [10:0] fifo_h2c_cmd_io_in_queue_io_upStream_bits_qid; // @[RegSlices.scala 64:35]
  wire  fifo_h2c_cmd_io_in_queue_io_upStream_bits_error; // @[RegSlices.scala 64:35]
  wire [7:0] fifo_h2c_cmd_io_in_queue_io_upStream_bits_func; // @[RegSlices.scala 64:35]
  wire [15:0] fifo_h2c_cmd_io_in_queue_io_upStream_bits_cidx; // @[RegSlices.scala 64:35]
  wire [2:0] fifo_h2c_cmd_io_in_queue_io_upStream_bits_port_id; // @[RegSlices.scala 64:35]
  wire  fifo_h2c_cmd_io_in_queue_io_upStream_bits_no_dma; // @[RegSlices.scala 64:35]
  wire  fifo_h2c_cmd_io_in_queue_io_downStream_ready; // @[RegSlices.scala 64:35]
  wire  fifo_h2c_cmd_io_in_queue_io_downStream_valid; // @[RegSlices.scala 64:35]
  wire [63:0] fifo_h2c_cmd_io_in_queue_io_downStream_bits_addr; // @[RegSlices.scala 64:35]
  wire [31:0] fifo_h2c_cmd_io_in_queue_io_downStream_bits_len; // @[RegSlices.scala 64:35]
  wire  fifo_h2c_cmd_io_in_queue_io_downStream_bits_eop; // @[RegSlices.scala 64:35]
  wire  fifo_h2c_cmd_io_in_queue_io_downStream_bits_sop; // @[RegSlices.scala 64:35]
  wire  fifo_h2c_cmd_io_in_queue_io_downStream_bits_mrkr_req; // @[RegSlices.scala 64:35]
  wire  fifo_h2c_cmd_io_in_queue_io_downStream_bits_sdi; // @[RegSlices.scala 64:35]
  wire [10:0] fifo_h2c_cmd_io_in_queue_io_downStream_bits_qid; // @[RegSlices.scala 64:35]
  wire  fifo_h2c_cmd_io_in_queue_io_downStream_bits_error; // @[RegSlices.scala 64:35]
  wire [7:0] fifo_h2c_cmd_io_in_queue_io_downStream_bits_func; // @[RegSlices.scala 64:35]
  wire [15:0] fifo_h2c_cmd_io_in_queue_io_downStream_bits_cidx; // @[RegSlices.scala 64:35]
  wire [2:0] fifo_h2c_cmd_io_in_queue_io_downStream_bits_port_id; // @[RegSlices.scala 64:35]
  wire  fifo_h2c_cmd_io_in_queue_io_downStream_bits_no_dma; // @[RegSlices.scala 64:35]
  wire  axil2reg_clock; // @[QDMADynamic.scala 86:76]
  wire  axil2reg_reset; // @[QDMADynamic.scala 86:76]
  wire  axil2reg_io_axi_aw_ready; // @[QDMADynamic.scala 86:76]
  wire  axil2reg_io_axi_aw_valid; // @[QDMADynamic.scala 86:76]
  wire [31:0] axil2reg_io_axi_aw_bits_addr; // @[QDMADynamic.scala 86:76]
  wire  axil2reg_io_axi_ar_ready; // @[QDMADynamic.scala 86:76]
  wire  axil2reg_io_axi_ar_valid; // @[QDMADynamic.scala 86:76]
  wire [31:0] axil2reg_io_axi_ar_bits_addr; // @[QDMADynamic.scala 86:76]
  wire  axil2reg_io_axi_w_ready; // @[QDMADynamic.scala 86:76]
  wire  axil2reg_io_axi_w_valid; // @[QDMADynamic.scala 86:76]
  wire [31:0] axil2reg_io_axi_w_bits_data; // @[QDMADynamic.scala 86:76]
  wire  axil2reg_io_axi_r_ready; // @[QDMADynamic.scala 86:76]
  wire  axil2reg_io_axi_r_valid; // @[QDMADynamic.scala 86:76]
  wire [31:0] axil2reg_io_axi_r_bits_data; // @[QDMADynamic.scala 86:76]
  wire [31:0] axil2reg_io_reg_control_0; // @[QDMADynamic.scala 86:76]
  wire [31:0] axil2reg_io_reg_control_8; // @[QDMADynamic.scala 86:76]
  wire [31:0] axil2reg_io_reg_control_9; // @[QDMADynamic.scala 86:76]
  wire [31:0] axil2reg_io_reg_control_10; // @[QDMADynamic.scala 86:76]
  wire [31:0] axil2reg_io_reg_control_11; // @[QDMADynamic.scala 86:76]
  wire [31:0] axil2reg_io_reg_control_12; // @[QDMADynamic.scala 86:76]
  wire [31:0] axil2reg_io_reg_control_13; // @[QDMADynamic.scala 86:76]
  wire [31:0] axil2reg_io_reg_control_14; // @[QDMADynamic.scala 86:76]
  wire [31:0] axil2reg_io_reg_status_300; // @[QDMADynamic.scala 86:76]
  wire [31:0] axil2reg_io_reg_status_400; // @[QDMADynamic.scala 86:76]
  wire [31:0] axil2reg_io_reg_status_401; // @[QDMADynamic.scala 86:76]
  wire [31:0] axil2reg_io_reg_status_402; // @[QDMADynamic.scala 86:76]
  wire [31:0] axil2reg_io_reg_status_403; // @[QDMADynamic.scala 86:76]
  wire [31:0] axil2reg_io_reg_status_404; // @[QDMADynamic.scala 86:76]
  wire [31:0] axil2reg_io_reg_status_405; // @[QDMADynamic.scala 86:76]
  wire [31:0] axil2reg_io_reg_status_406; // @[QDMADynamic.scala 86:76]
  wire [31:0] axil2reg_io_reg_status_407; // @[QDMADynamic.scala 86:76]
  wire [31:0] axil2reg_io_reg_status_408; // @[QDMADynamic.scala 86:76]
  wire [31:0] axil2reg_io_reg_status_409; // @[QDMADynamic.scala 86:76]
  wire [31:0] axil2reg_io_reg_status_410; // @[QDMADynamic.scala 86:76]
  wire [31:0] axil2reg_io_reg_status_411; // @[QDMADynamic.scala 86:76]
  wire [31:0] axil2reg_io_reg_status_412; // @[QDMADynamic.scala 86:76]
  wire [31:0] axil2reg_io_reg_status_413; // @[QDMADynamic.scala 86:76]
  wire [31:0] axil2reg_io_reg_status_414; // @[QDMADynamic.scala 86:76]
  wire  io_axib_cvt_aw_io_in_clk; // @[XConverter.scala 61:33]
  wire  io_axib_cvt_aw_io_out_clk; // @[XConverter.scala 61:33]
  wire  io_axib_cvt_aw_io_rstn; // @[XConverter.scala 61:33]
  wire  io_axib_cvt_aw_io_in_ready; // @[XConverter.scala 61:33]
  wire  io_axib_cvt_aw_io_in_valid; // @[XConverter.scala 61:33]
  wire [63:0] io_axib_cvt_aw_io_in_bits_addr; // @[XConverter.scala 61:33]
  wire [1:0] io_axib_cvt_aw_io_in_bits_burst; // @[XConverter.scala 61:33]
  wire [3:0] io_axib_cvt_aw_io_in_bits_cache; // @[XConverter.scala 61:33]
  wire [3:0] io_axib_cvt_aw_io_in_bits_id; // @[XConverter.scala 61:33]
  wire [7:0] io_axib_cvt_aw_io_in_bits_len; // @[XConverter.scala 61:33]
  wire  io_axib_cvt_aw_io_in_bits_lock; // @[XConverter.scala 61:33]
  wire [2:0] io_axib_cvt_aw_io_in_bits_prot; // @[XConverter.scala 61:33]
  wire [2:0] io_axib_cvt_aw_io_in_bits_size; // @[XConverter.scala 61:33]
  wire  io_axib_cvt_aw_io_out_ready; // @[XConverter.scala 61:33]
  wire  io_axib_cvt_aw_io_out_valid; // @[XConverter.scala 61:33]
  wire [63:0] io_axib_cvt_aw_io_out_bits_addr; // @[XConverter.scala 61:33]
  wire  io_axib_cvt_ar_io_in_clk; // @[XConverter.scala 61:33]
  wire  io_axib_cvt_ar_io_out_clk; // @[XConverter.scala 61:33]
  wire  io_axib_cvt_ar_io_rstn; // @[XConverter.scala 61:33]
  wire  io_axib_cvt_ar_io_in_ready; // @[XConverter.scala 61:33]
  wire  io_axib_cvt_ar_io_in_valid; // @[XConverter.scala 61:33]
  wire [63:0] io_axib_cvt_ar_io_in_bits_addr; // @[XConverter.scala 61:33]
  wire [1:0] io_axib_cvt_ar_io_in_bits_burst; // @[XConverter.scala 61:33]
  wire [3:0] io_axib_cvt_ar_io_in_bits_cache; // @[XConverter.scala 61:33]
  wire [3:0] io_axib_cvt_ar_io_in_bits_id; // @[XConverter.scala 61:33]
  wire [7:0] io_axib_cvt_ar_io_in_bits_len; // @[XConverter.scala 61:33]
  wire  io_axib_cvt_ar_io_in_bits_lock; // @[XConverter.scala 61:33]
  wire [2:0] io_axib_cvt_ar_io_in_bits_prot; // @[XConverter.scala 61:33]
  wire [2:0] io_axib_cvt_ar_io_in_bits_size; // @[XConverter.scala 61:33]
  wire  io_axib_cvt_ar_io_out_ready; // @[XConverter.scala 61:33]
  wire  io_axib_cvt_ar_io_out_valid; // @[XConverter.scala 61:33]
  wire [63:0] io_axib_cvt_ar_io_out_bits_addr; // @[XConverter.scala 61:33]
  wire  io_axib_cvt_w_io_in_clk; // @[XConverter.scala 61:33]
  wire  io_axib_cvt_w_io_out_clk; // @[XConverter.scala 61:33]
  wire  io_axib_cvt_w_io_rstn; // @[XConverter.scala 61:33]
  wire  io_axib_cvt_w_io_in_ready; // @[XConverter.scala 61:33]
  wire  io_axib_cvt_w_io_in_valid; // @[XConverter.scala 61:33]
  wire [511:0] io_axib_cvt_w_io_in_bits_data; // @[XConverter.scala 61:33]
  wire  io_axib_cvt_w_io_in_bits_last; // @[XConverter.scala 61:33]
  wire [63:0] io_axib_cvt_w_io_in_bits_strb; // @[XConverter.scala 61:33]
  wire  io_axib_cvt_w_io_out_ready; // @[XConverter.scala 61:33]
  wire  io_axib_cvt_w_io_out_valid; // @[XConverter.scala 61:33]
  wire [511:0] io_axib_cvt_w_io_out_bits_data; // @[XConverter.scala 61:33]
  wire  io_axib_cvt_r_io_in_clk; // @[XConverter.scala 61:33]
  wire  io_axib_cvt_r_io_out_clk; // @[XConverter.scala 61:33]
  wire  io_axib_cvt_r_io_rstn; // @[XConverter.scala 61:33]
  wire  io_axib_cvt_r_io_in_ready; // @[XConverter.scala 61:33]
  wire [511:0] io_axib_cvt_r_io_in_bits_data; // @[XConverter.scala 61:33]
  wire  io_axib_cvt_r_io_out_ready; // @[XConverter.scala 61:33]
  wire  io_axib_cvt_r_io_out_valid; // @[XConverter.scala 61:33]
  wire [511:0] io_axib_cvt_r_io_out_bits_data; // @[XConverter.scala 61:33]
  wire  io_axib_cvt_r_io_out_bits_last; // @[XConverter.scala 61:33]
  wire [1:0] io_axib_cvt_r_io_out_bits_resp; // @[XConverter.scala 61:33]
  wire [3:0] io_axib_cvt_r_io_out_bits_id; // @[XConverter.scala 61:33]
  wire  io_axib_cvt_b_io_in_clk; // @[XConverter.scala 61:33]
  wire  io_axib_cvt_b_io_out_clk; // @[XConverter.scala 61:33]
  wire  io_axib_cvt_b_io_rstn; // @[XConverter.scala 61:33]
  wire  io_axib_cvt_b_io_out_ready; // @[XConverter.scala 61:33]
  wire  io_axib_cvt_b_io_out_valid; // @[XConverter.scala 61:33]
  wire [3:0] io_axib_cvt_b_io_out_bits_id; // @[XConverter.scala 61:33]
  wire [1:0] io_axib_cvt_b_io_out_bits_resp; // @[XConverter.scala 61:33]
  wire  axil2reg_io_axi_cvt_aw_io_in_clk; // @[XConverter.scala 61:33]
  wire  axil2reg_io_axi_cvt_aw_io_out_clk; // @[XConverter.scala 61:33]
  wire  axil2reg_io_axi_cvt_aw_io_rstn; // @[XConverter.scala 61:33]
  wire  axil2reg_io_axi_cvt_aw_io_in_ready; // @[XConverter.scala 61:33]
  wire  axil2reg_io_axi_cvt_aw_io_in_valid; // @[XConverter.scala 61:33]
  wire [31:0] axil2reg_io_axi_cvt_aw_io_in_bits_addr; // @[XConverter.scala 61:33]
  wire  axil2reg_io_axi_cvt_aw_io_out_ready; // @[XConverter.scala 61:33]
  wire  axil2reg_io_axi_cvt_aw_io_out_valid; // @[XConverter.scala 61:33]
  wire [31:0] axil2reg_io_axi_cvt_aw_io_out_bits_addr; // @[XConverter.scala 61:33]
  wire  axil2reg_io_axi_cvt_ar_io_in_clk; // @[XConverter.scala 61:33]
  wire  axil2reg_io_axi_cvt_ar_io_out_clk; // @[XConverter.scala 61:33]
  wire  axil2reg_io_axi_cvt_ar_io_rstn; // @[XConverter.scala 61:33]
  wire  axil2reg_io_axi_cvt_ar_io_in_ready; // @[XConverter.scala 61:33]
  wire  axil2reg_io_axi_cvt_ar_io_in_valid; // @[XConverter.scala 61:33]
  wire [31:0] axil2reg_io_axi_cvt_ar_io_in_bits_addr; // @[XConverter.scala 61:33]
  wire  axil2reg_io_axi_cvt_ar_io_out_ready; // @[XConverter.scala 61:33]
  wire  axil2reg_io_axi_cvt_ar_io_out_valid; // @[XConverter.scala 61:33]
  wire [31:0] axil2reg_io_axi_cvt_ar_io_out_bits_addr; // @[XConverter.scala 61:33]
  wire  axil2reg_io_axi_cvt_w_io_in_clk; // @[XConverter.scala 61:33]
  wire  axil2reg_io_axi_cvt_w_io_out_clk; // @[XConverter.scala 61:33]
  wire  axil2reg_io_axi_cvt_w_io_rstn; // @[XConverter.scala 61:33]
  wire  axil2reg_io_axi_cvt_w_io_in_ready; // @[XConverter.scala 61:33]
  wire  axil2reg_io_axi_cvt_w_io_in_valid; // @[XConverter.scala 61:33]
  wire [31:0] axil2reg_io_axi_cvt_w_io_in_bits_data; // @[XConverter.scala 61:33]
  wire [3:0] axil2reg_io_axi_cvt_w_io_in_bits_strb; // @[XConverter.scala 61:33]
  wire  axil2reg_io_axi_cvt_w_io_out_ready; // @[XConverter.scala 61:33]
  wire  axil2reg_io_axi_cvt_w_io_out_valid; // @[XConverter.scala 61:33]
  wire [31:0] axil2reg_io_axi_cvt_w_io_out_bits_data; // @[XConverter.scala 61:33]
  wire  axil2reg_io_axi_cvt_r_io_in_clk; // @[XConverter.scala 61:33]
  wire  axil2reg_io_axi_cvt_r_io_out_clk; // @[XConverter.scala 61:33]
  wire  axil2reg_io_axi_cvt_r_io_rstn; // @[XConverter.scala 61:33]
  wire  axil2reg_io_axi_cvt_r_io_in_ready; // @[XConverter.scala 61:33]
  wire  axil2reg_io_axi_cvt_r_io_in_valid; // @[XConverter.scala 61:33]
  wire [31:0] axil2reg_io_axi_cvt_r_io_in_bits_data; // @[XConverter.scala 61:33]
  wire  axil2reg_io_axi_cvt_r_io_out_ready; // @[XConverter.scala 61:33]
  wire  axil2reg_io_axi_cvt_r_io_out_valid; // @[XConverter.scala 61:33]
  wire [31:0] axil2reg_io_axi_cvt_r_io_out_bits_data; // @[XConverter.scala 61:33]
  wire [1:0] axil2reg_io_axi_cvt_r_io_out_bits_resp; // @[XConverter.scala 61:33]
  wire  axil2reg_io_axi_cvt_b_io_in_clk; // @[XConverter.scala 61:33]
  wire  axil2reg_io_axi_cvt_b_io_out_clk; // @[XConverter.scala 61:33]
  wire  axil2reg_io_axi_cvt_b_io_rstn; // @[XConverter.scala 61:33]
  wire  axil2reg_io_axi_cvt_b_io_out_ready; // @[XConverter.scala 61:33]
  wire  axil2reg_io_axi_cvt_b_io_out_valid; // @[XConverter.scala 61:33]
  wire [1:0] axil2reg_io_axi_cvt_b_io_out_bits_resp; // @[XConverter.scala 61:33]
  wire  boundary_split_clock; // @[QDMADynamic.scala 116:82]
  wire  boundary_split_reset; // @[QDMADynamic.scala 116:82]
  wire  boundary_split_io_cmd_in_ready; // @[QDMADynamic.scala 116:82]
  wire  boundary_split_io_cmd_in_valid; // @[QDMADynamic.scala 116:82]
  wire [63:0] boundary_split_io_cmd_in_bits_addr; // @[QDMADynamic.scala 116:82]
  wire [10:0] boundary_split_io_cmd_in_bits_qid; // @[QDMADynamic.scala 116:82]
  wire  boundary_split_io_cmd_in_bits_error; // @[QDMADynamic.scala 116:82]
  wire [7:0] boundary_split_io_cmd_in_bits_func; // @[QDMADynamic.scala 116:82]
  wire [2:0] boundary_split_io_cmd_in_bits_port_id; // @[QDMADynamic.scala 116:82]
  wire [6:0] boundary_split_io_cmd_in_bits_pfch_tag; // @[QDMADynamic.scala 116:82]
  wire [31:0] boundary_split_io_cmd_in_bits_len; // @[QDMADynamic.scala 116:82]
  wire  boundary_split_io_data_out_ready; // @[QDMADynamic.scala 116:82]
  wire  boundary_split_io_data_out_valid; // @[QDMADynamic.scala 116:82]
  wire [511:0] boundary_split_io_data_out_bits_data; // @[QDMADynamic.scala 116:82]
  wire [31:0] boundary_split_io_data_out_bits_tcrc; // @[QDMADynamic.scala 116:82]
  wire  boundary_split_io_data_out_bits_ctrl_marker; // @[QDMADynamic.scala 116:82]
  wire [6:0] boundary_split_io_data_out_bits_ctrl_ecc; // @[QDMADynamic.scala 116:82]
  wire [31:0] boundary_split_io_data_out_bits_ctrl_len; // @[QDMADynamic.scala 116:82]
  wire [2:0] boundary_split_io_data_out_bits_ctrl_port_id; // @[QDMADynamic.scala 116:82]
  wire [10:0] boundary_split_io_data_out_bits_ctrl_qid; // @[QDMADynamic.scala 116:82]
  wire  boundary_split_io_data_out_bits_ctrl_has_cmpt; // @[QDMADynamic.scala 116:82]
  wire  boundary_split_io_data_out_bits_last; // @[QDMADynamic.scala 116:82]
  wire [5:0] boundary_split_io_data_out_bits_mty; // @[QDMADynamic.scala 116:82]
  wire  boundary_split_io_cmd_out_ready; // @[QDMADynamic.scala 116:82]
  wire  boundary_split_io_cmd_out_valid; // @[QDMADynamic.scala 116:82]
  wire [63:0] boundary_split_io_cmd_out_bits_addr; // @[QDMADynamic.scala 116:82]
  wire [10:0] boundary_split_io_cmd_out_bits_qid; // @[QDMADynamic.scala 116:82]
  wire  boundary_split_io_cmd_out_bits_error; // @[QDMADynamic.scala 116:82]
  wire [7:0] boundary_split_io_cmd_out_bits_func; // @[QDMADynamic.scala 116:82]
  wire [2:0] boundary_split_io_cmd_out_bits_port_id; // @[QDMADynamic.scala 116:82]
  wire [6:0] boundary_split_io_cmd_out_bits_pfch_tag; // @[QDMADynamic.scala 116:82]
  wire [31:0] boundary_split_io_cmd_out_bits_len; // @[QDMADynamic.scala 116:82]
  wire  _fifo_h2c_data_io_in_T = ~io_qdma_port_axi_aresetn; // @[QDMADynamic.scala 52:73]
  wire  _T = ~io_user_arstn; // @[QDMADynamic.scala 62:73]
  reg  wr_tlb_valid_REG; // @[QDMADynamic.scala 81:99]
  reg  wr_tlb_valid_REG_1; // @[QDMADynamic.scala 81:90]
  wire  _T_6 = _T | sw_reset_pad_O; // @[QDMADynamic.scala 122:55]
  reg [31:0] counter; // @[Collector.scala 169:42]
  reg [31:0] counter_1; // @[Collector.scala 169:42]
  wire  _T_8 = io_h2c_cmd_ready & io_h2c_cmd_valid; // @[Decoupled.scala 40:37]
  wire [31:0] _counter_T_3 = counter_1 + 32'h1; // @[Collector.scala 171:51]
  reg [31:0] counter_2; // @[Collector.scala 169:42]
  reg [31:0] counter_3; // @[Collector.scala 169:42]
  wire [31:0] _counter_T_7 = counter_3 + 32'h1; // @[Collector.scala 171:51]
  wire  _T_12 = _fifo_h2c_data_io_in_T | sw_reset_pad_O; // @[QDMADynamic.scala 129:49]
  reg [31:0] counter_4; // @[Collector.scala 169:42]
  wire  _T_13 = fifo_c2h_cmd_io_out_ready & fifo_c2h_cmd_io_out_valid; // @[Decoupled.scala 40:37]
  wire [31:0] _counter_T_9 = counter_4 + 32'h1; // @[Collector.scala 171:51]
  reg [31:0] counter_5; // @[Collector.scala 169:42]
  wire  _T_14 = fifo_h2c_cmd_io__out_ready & fifo_h2c_cmd_io__out_valid; // @[Decoupled.scala 40:37]
  wire [31:0] _counter_T_11 = counter_5 + 32'h1; // @[Collector.scala 171:51]
  reg [31:0] counter_6; // @[Collector.scala 169:42]
  wire  _T_15 = fifo_c2h_data_io__out_ready & fifo_c2h_data_io__out_valid; // @[Decoupled.scala 40:37]
  wire [31:0] _counter_T_13 = counter_6 + 32'h1; // @[Collector.scala 171:51]
  reg [31:0] counter_7; // @[Collector.scala 169:42]
  wire  _T_16 = fifo_h2c_data_io__in_ready & fifo_h2c_data_io__in_valid; // @[Decoupled.scala 40:37]
  wire [31:0] _counter_T_15 = counter_7 + 32'h1; // @[Collector.scala 171:51]
  BUFG sw_reset_pad ( // @[Buf.scala 33:34]
    .O(sw_reset_pad_O),
    .I(sw_reset_pad_I)
  );
  XConverter fifo_h2c_data ( // @[XConverter.scala 61:33]
    .io__in_clk(fifo_h2c_data_io__in_clk),
    .io__out_clk(fifo_h2c_data_io__out_clk),
    .io__rstn(fifo_h2c_data_io__rstn),
    .io__in_ready(fifo_h2c_data_io__in_ready),
    .io__in_valid(fifo_h2c_data_io__in_valid),
    .io__in_bits_data(fifo_h2c_data_io__in_bits_data),
    .io__in_bits_tcrc(fifo_h2c_data_io__in_bits_tcrc),
    .io__in_bits_tuser_qid(fifo_h2c_data_io__in_bits_tuser_qid),
    .io__in_bits_tuser_port_id(fifo_h2c_data_io__in_bits_tuser_port_id),
    .io__in_bits_tuser_err(fifo_h2c_data_io__in_bits_tuser_err),
    .io__in_bits_tuser_mdata(fifo_h2c_data_io__in_bits_tuser_mdata),
    .io__in_bits_tuser_mty(fifo_h2c_data_io__in_bits_tuser_mty),
    .io__in_bits_tuser_zero_byte(fifo_h2c_data_io__in_bits_tuser_zero_byte),
    .io__in_bits_last(fifo_h2c_data_io__in_bits_last),
    .io__out_valid(fifo_h2c_data_io__out_valid),
    .io_in_ready(fifo_h2c_data_io_in_ready),
    .io_in_valid(fifo_h2c_data_io_in_valid)
  );
  RegSlice fifo_h2c_data_io_in_queue ( // @[RegSlices.scala 64:35]
    .clock(fifo_h2c_data_io_in_queue_clock),
    .reset(fifo_h2c_data_io_in_queue_reset),
    .io_upStream_ready(fifo_h2c_data_io_in_queue_io_upStream_ready),
    .io_upStream_valid(fifo_h2c_data_io_in_queue_io_upStream_valid),
    .io_upStream_bits_data(fifo_h2c_data_io_in_queue_io_upStream_bits_data),
    .io_upStream_bits_tcrc(fifo_h2c_data_io_in_queue_io_upStream_bits_tcrc),
    .io_upStream_bits_tuser_qid(fifo_h2c_data_io_in_queue_io_upStream_bits_tuser_qid),
    .io_upStream_bits_tuser_port_id(fifo_h2c_data_io_in_queue_io_upStream_bits_tuser_port_id),
    .io_upStream_bits_tuser_err(fifo_h2c_data_io_in_queue_io_upStream_bits_tuser_err),
    .io_upStream_bits_tuser_mdata(fifo_h2c_data_io_in_queue_io_upStream_bits_tuser_mdata),
    .io_upStream_bits_tuser_mty(fifo_h2c_data_io_in_queue_io_upStream_bits_tuser_mty),
    .io_upStream_bits_tuser_zero_byte(fifo_h2c_data_io_in_queue_io_upStream_bits_tuser_zero_byte),
    .io_upStream_bits_last(fifo_h2c_data_io_in_queue_io_upStream_bits_last),
    .io_downStream_ready(fifo_h2c_data_io_in_queue_io_downStream_ready),
    .io_downStream_valid(fifo_h2c_data_io_in_queue_io_downStream_valid),
    .io_downStream_bits_data(fifo_h2c_data_io_in_queue_io_downStream_bits_data),
    .io_downStream_bits_tcrc(fifo_h2c_data_io_in_queue_io_downStream_bits_tcrc),
    .io_downStream_bits_tuser_qid(fifo_h2c_data_io_in_queue_io_downStream_bits_tuser_qid),
    .io_downStream_bits_tuser_port_id(fifo_h2c_data_io_in_queue_io_downStream_bits_tuser_port_id),
    .io_downStream_bits_tuser_err(fifo_h2c_data_io_in_queue_io_downStream_bits_tuser_err),
    .io_downStream_bits_tuser_mdata(fifo_h2c_data_io_in_queue_io_downStream_bits_tuser_mdata),
    .io_downStream_bits_tuser_mty(fifo_h2c_data_io_in_queue_io_downStream_bits_tuser_mty),
    .io_downStream_bits_tuser_zero_byte(fifo_h2c_data_io_in_queue_io_downStream_bits_tuser_zero_byte),
    .io_downStream_bits_last(fifo_h2c_data_io_in_queue_io_downStream_bits_last)
  );
  XConverter_1 fifo_c2h_data ( // @[XConverter.scala 61:33]
    .io__in_clk(fifo_c2h_data_io__in_clk),
    .io__out_clk(fifo_c2h_data_io__out_clk),
    .io__rstn(fifo_c2h_data_io__rstn),
    .io__in_ready(fifo_c2h_data_io__in_ready),
    .io__in_valid(fifo_c2h_data_io__in_valid),
    .io__in_bits_data(fifo_c2h_data_io__in_bits_data),
    .io__in_bits_tcrc(fifo_c2h_data_io__in_bits_tcrc),
    .io__in_bits_ctrl_marker(fifo_c2h_data_io__in_bits_ctrl_marker),
    .io__in_bits_ctrl_ecc(fifo_c2h_data_io__in_bits_ctrl_ecc),
    .io__in_bits_ctrl_len(fifo_c2h_data_io__in_bits_ctrl_len),
    .io__in_bits_ctrl_port_id(fifo_c2h_data_io__in_bits_ctrl_port_id),
    .io__in_bits_ctrl_qid(fifo_c2h_data_io__in_bits_ctrl_qid),
    .io__in_bits_ctrl_has_cmpt(fifo_c2h_data_io__in_bits_ctrl_has_cmpt),
    .io__in_bits_last(fifo_c2h_data_io__in_bits_last),
    .io__in_bits_mty(fifo_c2h_data_io__in_bits_mty),
    .io__out_ready(fifo_c2h_data_io__out_ready),
    .io__out_valid(fifo_c2h_data_io__out_valid),
    .io__out_bits_data(fifo_c2h_data_io__out_bits_data),
    .io__out_bits_tcrc(fifo_c2h_data_io__out_bits_tcrc),
    .io__out_bits_ctrl_marker(fifo_c2h_data_io__out_bits_ctrl_marker),
    .io__out_bits_ctrl_ecc(fifo_c2h_data_io__out_bits_ctrl_ecc),
    .io__out_bits_ctrl_len(fifo_c2h_data_io__out_bits_ctrl_len),
    .io__out_bits_ctrl_port_id(fifo_c2h_data_io__out_bits_ctrl_port_id),
    .io__out_bits_ctrl_qid(fifo_c2h_data_io__out_bits_ctrl_qid),
    .io__out_bits_ctrl_has_cmpt(fifo_c2h_data_io__out_bits_ctrl_has_cmpt),
    .io__out_bits_last(fifo_c2h_data_io__out_bits_last),
    .io__out_bits_mty(fifo_c2h_data_io__out_bits_mty),
    .io_out_ready(fifo_c2h_data_io_out_ready),
    .io_out_valid_0(fifo_c2h_data_io_out_valid_0)
  );
  RegSlice_1 fifo_c2h_data_out_queue ( // @[RegSlices.scala 64:35]
    .clock(fifo_c2h_data_out_queue_clock),
    .reset(fifo_c2h_data_out_queue_reset),
    .io_upStream_ready(fifo_c2h_data_out_queue_io_upStream_ready),
    .io_upStream_valid(fifo_c2h_data_out_queue_io_upStream_valid),
    .io_upStream_bits_data(fifo_c2h_data_out_queue_io_upStream_bits_data),
    .io_upStream_bits_tcrc(fifo_c2h_data_out_queue_io_upStream_bits_tcrc),
    .io_upStream_bits_ctrl_marker(fifo_c2h_data_out_queue_io_upStream_bits_ctrl_marker),
    .io_upStream_bits_ctrl_ecc(fifo_c2h_data_out_queue_io_upStream_bits_ctrl_ecc),
    .io_upStream_bits_ctrl_len(fifo_c2h_data_out_queue_io_upStream_bits_ctrl_len),
    .io_upStream_bits_ctrl_port_id(fifo_c2h_data_out_queue_io_upStream_bits_ctrl_port_id),
    .io_upStream_bits_ctrl_qid(fifo_c2h_data_out_queue_io_upStream_bits_ctrl_qid),
    .io_upStream_bits_ctrl_has_cmpt(fifo_c2h_data_out_queue_io_upStream_bits_ctrl_has_cmpt),
    .io_upStream_bits_last(fifo_c2h_data_out_queue_io_upStream_bits_last),
    .io_upStream_bits_mty(fifo_c2h_data_out_queue_io_upStream_bits_mty),
    .io_downStream_ready(fifo_c2h_data_out_queue_io_downStream_ready),
    .io_downStream_valid(fifo_c2h_data_out_queue_io_downStream_valid),
    .io_downStream_bits_data(fifo_c2h_data_out_queue_io_downStream_bits_data),
    .io_downStream_bits_tcrc(fifo_c2h_data_out_queue_io_downStream_bits_tcrc),
    .io_downStream_bits_ctrl_marker(fifo_c2h_data_out_queue_io_downStream_bits_ctrl_marker),
    .io_downStream_bits_ctrl_ecc(fifo_c2h_data_out_queue_io_downStream_bits_ctrl_ecc),
    .io_downStream_bits_ctrl_len(fifo_c2h_data_out_queue_io_downStream_bits_ctrl_len),
    .io_downStream_bits_ctrl_port_id(fifo_c2h_data_out_queue_io_downStream_bits_ctrl_port_id),
    .io_downStream_bits_ctrl_qid(fifo_c2h_data_out_queue_io_downStream_bits_ctrl_qid),
    .io_downStream_bits_ctrl_has_cmpt(fifo_c2h_data_out_queue_io_downStream_bits_ctrl_has_cmpt),
    .io_downStream_bits_last(fifo_c2h_data_out_queue_io_downStream_bits_last),
    .io_downStream_bits_mty(fifo_c2h_data_out_queue_io_downStream_bits_mty)
  );
  XConverter_2 fifo_h2c_cmd ( // @[XConverter.scala 61:33]
    .io__in_clk(fifo_h2c_cmd_io__in_clk),
    .io__out_clk(fifo_h2c_cmd_io__out_clk),
    .io__rstn(fifo_h2c_cmd_io__rstn),
    .io__in_ready(fifo_h2c_cmd_io__in_ready),
    .io__in_valid(fifo_h2c_cmd_io__in_valid),
    .io__in_bits_addr(fifo_h2c_cmd_io__in_bits_addr),
    .io__in_bits_len(fifo_h2c_cmd_io__in_bits_len),
    .io__in_bits_eop(fifo_h2c_cmd_io__in_bits_eop),
    .io__in_bits_sop(fifo_h2c_cmd_io__in_bits_sop),
    .io__in_bits_mrkr_req(fifo_h2c_cmd_io__in_bits_mrkr_req),
    .io__in_bits_sdi(fifo_h2c_cmd_io__in_bits_sdi),
    .io__in_bits_qid(fifo_h2c_cmd_io__in_bits_qid),
    .io__in_bits_error(fifo_h2c_cmd_io__in_bits_error),
    .io__in_bits_func(fifo_h2c_cmd_io__in_bits_func),
    .io__in_bits_cidx(fifo_h2c_cmd_io__in_bits_cidx),
    .io__in_bits_port_id(fifo_h2c_cmd_io__in_bits_port_id),
    .io__in_bits_no_dma(fifo_h2c_cmd_io__in_bits_no_dma),
    .io__out_ready(fifo_h2c_cmd_io__out_ready),
    .io__out_valid(fifo_h2c_cmd_io__out_valid),
    .io__out_bits_addr(fifo_h2c_cmd_io__out_bits_addr),
    .io__out_bits_len(fifo_h2c_cmd_io__out_bits_len),
    .io__out_bits_eop(fifo_h2c_cmd_io__out_bits_eop),
    .io__out_bits_sop(fifo_h2c_cmd_io__out_bits_sop),
    .io__out_bits_mrkr_req(fifo_h2c_cmd_io__out_bits_mrkr_req),
    .io__out_bits_sdi(fifo_h2c_cmd_io__out_bits_sdi),
    .io__out_bits_qid(fifo_h2c_cmd_io__out_bits_qid),
    .io__out_bits_error(fifo_h2c_cmd_io__out_bits_error),
    .io__out_bits_func(fifo_h2c_cmd_io__out_bits_func),
    .io__out_bits_cidx(fifo_h2c_cmd_io__out_bits_cidx),
    .io__out_bits_port_id(fifo_h2c_cmd_io__out_bits_port_id),
    .io__out_bits_no_dma(fifo_h2c_cmd_io__out_bits_no_dma),
    .io_out_valid(fifo_h2c_cmd_io_out_valid),
    .io_out_ready_1(fifo_h2c_cmd_io_out_ready_1)
  );
  RegSlice_2 fifo_h2c_cmd_out_queue ( // @[RegSlices.scala 64:35]
    .clock(fifo_h2c_cmd_out_queue_clock),
    .reset(fifo_h2c_cmd_out_queue_reset),
    .io_upStream_ready(fifo_h2c_cmd_out_queue_io_upStream_ready),
    .io_upStream_valid(fifo_h2c_cmd_out_queue_io_upStream_valid),
    .io_upStream_bits_addr(fifo_h2c_cmd_out_queue_io_upStream_bits_addr),
    .io_upStream_bits_len(fifo_h2c_cmd_out_queue_io_upStream_bits_len),
    .io_upStream_bits_eop(fifo_h2c_cmd_out_queue_io_upStream_bits_eop),
    .io_upStream_bits_sop(fifo_h2c_cmd_out_queue_io_upStream_bits_sop),
    .io_upStream_bits_mrkr_req(fifo_h2c_cmd_out_queue_io_upStream_bits_mrkr_req),
    .io_upStream_bits_sdi(fifo_h2c_cmd_out_queue_io_upStream_bits_sdi),
    .io_upStream_bits_qid(fifo_h2c_cmd_out_queue_io_upStream_bits_qid),
    .io_upStream_bits_error(fifo_h2c_cmd_out_queue_io_upStream_bits_error),
    .io_upStream_bits_func(fifo_h2c_cmd_out_queue_io_upStream_bits_func),
    .io_upStream_bits_cidx(fifo_h2c_cmd_out_queue_io_upStream_bits_cidx),
    .io_upStream_bits_port_id(fifo_h2c_cmd_out_queue_io_upStream_bits_port_id),
    .io_upStream_bits_no_dma(fifo_h2c_cmd_out_queue_io_upStream_bits_no_dma),
    .io_downStream_ready(fifo_h2c_cmd_out_queue_io_downStream_ready),
    .io_downStream_valid(fifo_h2c_cmd_out_queue_io_downStream_valid),
    .io_downStream_bits_addr(fifo_h2c_cmd_out_queue_io_downStream_bits_addr),
    .io_downStream_bits_len(fifo_h2c_cmd_out_queue_io_downStream_bits_len),
    .io_downStream_bits_eop(fifo_h2c_cmd_out_queue_io_downStream_bits_eop),
    .io_downStream_bits_sop(fifo_h2c_cmd_out_queue_io_downStream_bits_sop),
    .io_downStream_bits_mrkr_req(fifo_h2c_cmd_out_queue_io_downStream_bits_mrkr_req),
    .io_downStream_bits_sdi(fifo_h2c_cmd_out_queue_io_downStream_bits_sdi),
    .io_downStream_bits_qid(fifo_h2c_cmd_out_queue_io_downStream_bits_qid),
    .io_downStream_bits_error(fifo_h2c_cmd_out_queue_io_downStream_bits_error),
    .io_downStream_bits_func(fifo_h2c_cmd_out_queue_io_downStream_bits_func),
    .io_downStream_bits_cidx(fifo_h2c_cmd_out_queue_io_downStream_bits_cidx),
    .io_downStream_bits_port_id(fifo_h2c_cmd_out_queue_io_downStream_bits_port_id),
    .io_downStream_bits_no_dma(fifo_h2c_cmd_out_queue_io_downStream_bits_no_dma)
  );
  XConverter_3 fifo_c2h_cmd ( // @[XConverter.scala 61:33]
    .io_in_clk(fifo_c2h_cmd_io_in_clk),
    .io_out_clk(fifo_c2h_cmd_io_out_clk),
    .io_rstn(fifo_c2h_cmd_io_rstn),
    .io_in_ready(fifo_c2h_cmd_io_in_ready),
    .io_in_valid(fifo_c2h_cmd_io_in_valid),
    .io_in_bits_addr(fifo_c2h_cmd_io_in_bits_addr),
    .io_in_bits_qid(fifo_c2h_cmd_io_in_bits_qid),
    .io_in_bits_error(fifo_c2h_cmd_io_in_bits_error),
    .io_in_bits_func(fifo_c2h_cmd_io_in_bits_func),
    .io_in_bits_port_id(fifo_c2h_cmd_io_in_bits_port_id),
    .io_in_bits_pfch_tag(fifo_c2h_cmd_io_in_bits_pfch_tag),
    .io_in_bits_len(fifo_c2h_cmd_io_in_bits_len),
    .io_out_ready(fifo_c2h_cmd_io_out_ready),
    .io_out_valid(fifo_c2h_cmd_io_out_valid),
    .io_out_bits_addr(fifo_c2h_cmd_io_out_bits_addr),
    .io_out_bits_qid(fifo_c2h_cmd_io_out_bits_qid),
    .io_out_bits_error(fifo_c2h_cmd_io_out_bits_error),
    .io_out_bits_func(fifo_c2h_cmd_io_out_bits_func),
    .io_out_bits_port_id(fifo_c2h_cmd_io_out_bits_port_id),
    .io_out_bits_pfch_tag(fifo_c2h_cmd_io_out_bits_pfch_tag),
    .io_out_bits_len(fifo_c2h_cmd_io_out_bits_len),
    .io_out_ready_0(fifo_c2h_cmd_io_out_ready_0),
    .io_out_valid_1(fifo_c2h_cmd_io_out_valid_1)
  );
  RegSlice_3 fifo_c2h_cmd_out_queue ( // @[RegSlices.scala 64:35]
    .clock(fifo_c2h_cmd_out_queue_clock),
    .reset(fifo_c2h_cmd_out_queue_reset),
    .io_upStream_ready(fifo_c2h_cmd_out_queue_io_upStream_ready),
    .io_upStream_valid(fifo_c2h_cmd_out_queue_io_upStream_valid),
    .io_upStream_bits_addr(fifo_c2h_cmd_out_queue_io_upStream_bits_addr),
    .io_upStream_bits_qid(fifo_c2h_cmd_out_queue_io_upStream_bits_qid),
    .io_upStream_bits_error(fifo_c2h_cmd_out_queue_io_upStream_bits_error),
    .io_upStream_bits_func(fifo_c2h_cmd_out_queue_io_upStream_bits_func),
    .io_upStream_bits_port_id(fifo_c2h_cmd_out_queue_io_upStream_bits_port_id),
    .io_upStream_bits_pfch_tag(fifo_c2h_cmd_out_queue_io_upStream_bits_pfch_tag),
    .io_upStream_bits_len(fifo_c2h_cmd_out_queue_io_upStream_bits_len),
    .io_downStream_ready(fifo_c2h_cmd_out_queue_io_downStream_ready),
    .io_downStream_valid(fifo_c2h_cmd_out_queue_io_downStream_valid),
    .io_downStream_bits_addr(fifo_c2h_cmd_out_queue_io_downStream_bits_addr),
    .io_downStream_bits_qid(fifo_c2h_cmd_out_queue_io_downStream_bits_qid),
    .io_downStream_bits_error(fifo_c2h_cmd_out_queue_io_downStream_bits_error),
    .io_downStream_bits_func(fifo_c2h_cmd_out_queue_io_downStream_bits_func),
    .io_downStream_bits_port_id(fifo_c2h_cmd_out_queue_io_downStream_bits_port_id),
    .io_downStream_bits_pfch_tag(fifo_c2h_cmd_out_queue_io_downStream_bits_pfch_tag),
    .io_downStream_bits_len(fifo_c2h_cmd_out_queue_io_downStream_bits_len)
  );
  CMDBoundaryCheck check_c2h ( // @[QDMADynamic.scala 62:95]
    .clock(check_c2h_clock),
    .reset(check_c2h_reset),
    .io_in_ready(check_c2h_io_in_ready),
    .io_in_valid(check_c2h_io_in_valid),
    .io_in_bits_addr(check_c2h_io_in_bits_addr),
    .io_in_bits_qid(check_c2h_io_in_bits_qid),
    .io_in_bits_error(check_c2h_io_in_bits_error),
    .io_in_bits_func(check_c2h_io_in_bits_func),
    .io_in_bits_port_id(check_c2h_io_in_bits_port_id),
    .io_in_bits_pfch_tag(check_c2h_io_in_bits_pfch_tag),
    .io_in_bits_len(check_c2h_io_in_bits_len),
    .io_out_ready(check_c2h_io_out_ready),
    .io_out_valid(check_c2h_io_out_valid),
    .io_out_bits_addr(check_c2h_io_out_bits_addr),
    .io_out_bits_qid(check_c2h_io_out_bits_qid),
    .io_out_bits_error(check_c2h_io_out_bits_error),
    .io_out_bits_func(check_c2h_io_out_bits_func),
    .io_out_bits_port_id(check_c2h_io_out_bits_port_id),
    .io_out_bits_pfch_tag(check_c2h_io_out_bits_pfch_tag),
    .io_out_bits_len(check_c2h_io_out_bits_len)
  );
  RegSlice_3 check_c2h_io_in_queue ( // @[RegSlices.scala 64:35]
    .clock(check_c2h_io_in_queue_clock),
    .reset(check_c2h_io_in_queue_reset),
    .io_upStream_ready(check_c2h_io_in_queue_io_upStream_ready),
    .io_upStream_valid(check_c2h_io_in_queue_io_upStream_valid),
    .io_upStream_bits_addr(check_c2h_io_in_queue_io_upStream_bits_addr),
    .io_upStream_bits_qid(check_c2h_io_in_queue_io_upStream_bits_qid),
    .io_upStream_bits_error(check_c2h_io_in_queue_io_upStream_bits_error),
    .io_upStream_bits_func(check_c2h_io_in_queue_io_upStream_bits_func),
    .io_upStream_bits_port_id(check_c2h_io_in_queue_io_upStream_bits_port_id),
    .io_upStream_bits_pfch_tag(check_c2h_io_in_queue_io_upStream_bits_pfch_tag),
    .io_upStream_bits_len(check_c2h_io_in_queue_io_upStream_bits_len),
    .io_downStream_ready(check_c2h_io_in_queue_io_downStream_ready),
    .io_downStream_valid(check_c2h_io_in_queue_io_downStream_valid),
    .io_downStream_bits_addr(check_c2h_io_in_queue_io_downStream_bits_addr),
    .io_downStream_bits_qid(check_c2h_io_in_queue_io_downStream_bits_qid),
    .io_downStream_bits_error(check_c2h_io_in_queue_io_downStream_bits_error),
    .io_downStream_bits_func(check_c2h_io_in_queue_io_downStream_bits_func),
    .io_downStream_bits_port_id(check_c2h_io_in_queue_io_downStream_bits_port_id),
    .io_downStream_bits_pfch_tag(check_c2h_io_in_queue_io_downStream_bits_pfch_tag),
    .io_downStream_bits_len(check_c2h_io_in_queue_io_downStream_bits_len)
  );
  CMDBoundaryCheck_1 check_h2c ( // @[QDMADynamic.scala 64:95]
    .clock(check_h2c_clock),
    .reset(check_h2c_reset),
    .io_in_ready(check_h2c_io_in_ready),
    .io_in_valid(check_h2c_io_in_valid),
    .io_in_bits_addr(check_h2c_io_in_bits_addr),
    .io_in_bits_len(check_h2c_io_in_bits_len),
    .io_in_bits_eop(check_h2c_io_in_bits_eop),
    .io_in_bits_sop(check_h2c_io_in_bits_sop),
    .io_in_bits_mrkr_req(check_h2c_io_in_bits_mrkr_req),
    .io_in_bits_sdi(check_h2c_io_in_bits_sdi),
    .io_in_bits_qid(check_h2c_io_in_bits_qid),
    .io_in_bits_error(check_h2c_io_in_bits_error),
    .io_in_bits_func(check_h2c_io_in_bits_func),
    .io_in_bits_cidx(check_h2c_io_in_bits_cidx),
    .io_in_bits_port_id(check_h2c_io_in_bits_port_id),
    .io_in_bits_no_dma(check_h2c_io_in_bits_no_dma),
    .io_out_ready(check_h2c_io_out_ready),
    .io_out_valid(check_h2c_io_out_valid),
    .io_out_bits_addr(check_h2c_io_out_bits_addr),
    .io_out_bits_len(check_h2c_io_out_bits_len),
    .io_out_bits_eop(check_h2c_io_out_bits_eop),
    .io_out_bits_sop(check_h2c_io_out_bits_sop),
    .io_out_bits_mrkr_req(check_h2c_io_out_bits_mrkr_req),
    .io_out_bits_sdi(check_h2c_io_out_bits_sdi),
    .io_out_bits_qid(check_h2c_io_out_bits_qid),
    .io_out_bits_error(check_h2c_io_out_bits_error),
    .io_out_bits_func(check_h2c_io_out_bits_func),
    .io_out_bits_cidx(check_h2c_io_out_bits_cidx),
    .io_out_bits_port_id(check_h2c_io_out_bits_port_id),
    .io_out_bits_no_dma(check_h2c_io_out_bits_no_dma)
  );
  RegSlice_2 check_h2c_io_in_queue ( // @[RegSlices.scala 64:35]
    .clock(check_h2c_io_in_queue_clock),
    .reset(check_h2c_io_in_queue_reset),
    .io_upStream_ready(check_h2c_io_in_queue_io_upStream_ready),
    .io_upStream_valid(check_h2c_io_in_queue_io_upStream_valid),
    .io_upStream_bits_addr(check_h2c_io_in_queue_io_upStream_bits_addr),
    .io_upStream_bits_len(check_h2c_io_in_queue_io_upStream_bits_len),
    .io_upStream_bits_eop(check_h2c_io_in_queue_io_upStream_bits_eop),
    .io_upStream_bits_sop(check_h2c_io_in_queue_io_upStream_bits_sop),
    .io_upStream_bits_mrkr_req(check_h2c_io_in_queue_io_upStream_bits_mrkr_req),
    .io_upStream_bits_sdi(check_h2c_io_in_queue_io_upStream_bits_sdi),
    .io_upStream_bits_qid(check_h2c_io_in_queue_io_upStream_bits_qid),
    .io_upStream_bits_error(check_h2c_io_in_queue_io_upStream_bits_error),
    .io_upStream_bits_func(check_h2c_io_in_queue_io_upStream_bits_func),
    .io_upStream_bits_cidx(check_h2c_io_in_queue_io_upStream_bits_cidx),
    .io_upStream_bits_port_id(check_h2c_io_in_queue_io_upStream_bits_port_id),
    .io_upStream_bits_no_dma(check_h2c_io_in_queue_io_upStream_bits_no_dma),
    .io_downStream_ready(check_h2c_io_in_queue_io_downStream_ready),
    .io_downStream_valid(check_h2c_io_in_queue_io_downStream_valid),
    .io_downStream_bits_addr(check_h2c_io_in_queue_io_downStream_bits_addr),
    .io_downStream_bits_len(check_h2c_io_in_queue_io_downStream_bits_len),
    .io_downStream_bits_eop(check_h2c_io_in_queue_io_downStream_bits_eop),
    .io_downStream_bits_sop(check_h2c_io_in_queue_io_downStream_bits_sop),
    .io_downStream_bits_mrkr_req(check_h2c_io_in_queue_io_downStream_bits_mrkr_req),
    .io_downStream_bits_sdi(check_h2c_io_in_queue_io_downStream_bits_sdi),
    .io_downStream_bits_qid(check_h2c_io_in_queue_io_downStream_bits_qid),
    .io_downStream_bits_error(check_h2c_io_in_queue_io_downStream_bits_error),
    .io_downStream_bits_func(check_h2c_io_in_queue_io_downStream_bits_func),
    .io_downStream_bits_cidx(check_h2c_io_in_queue_io_downStream_bits_cidx),
    .io_downStream_bits_port_id(check_h2c_io_in_queue_io_downStream_bits_port_id),
    .io_downStream_bits_no_dma(check_h2c_io_in_queue_io_downStream_bits_no_dma)
  );
  TLB tlb ( // @[QDMADynamic.scala 67:71]
    .clock(tlb_clock),
    .reset(tlb_reset),
    .io__wr_tlb_ready(tlb_io__wr_tlb_ready),
    .io__wr_tlb_valid(tlb_io__wr_tlb_valid),
    .io__wr_tlb_bits_vaddr_high(tlb_io__wr_tlb_bits_vaddr_high),
    .io__wr_tlb_bits_vaddr_low(tlb_io__wr_tlb_bits_vaddr_low),
    .io__wr_tlb_bits_paddr_high(tlb_io__wr_tlb_bits_paddr_high),
    .io__wr_tlb_bits_paddr_low(tlb_io__wr_tlb_bits_paddr_low),
    .io__wr_tlb_bits_is_base(tlb_io__wr_tlb_bits_is_base),
    .io__h2c_in_ready(tlb_io__h2c_in_ready),
    .io__h2c_in_valid(tlb_io__h2c_in_valid),
    .io__h2c_in_bits_addr(tlb_io__h2c_in_bits_addr),
    .io__h2c_in_bits_len(tlb_io__h2c_in_bits_len),
    .io__h2c_in_bits_eop(tlb_io__h2c_in_bits_eop),
    .io__h2c_in_bits_sop(tlb_io__h2c_in_bits_sop),
    .io__h2c_in_bits_mrkr_req(tlb_io__h2c_in_bits_mrkr_req),
    .io__h2c_in_bits_sdi(tlb_io__h2c_in_bits_sdi),
    .io__h2c_in_bits_qid(tlb_io__h2c_in_bits_qid),
    .io__h2c_in_bits_error(tlb_io__h2c_in_bits_error),
    .io__h2c_in_bits_func(tlb_io__h2c_in_bits_func),
    .io__h2c_in_bits_cidx(tlb_io__h2c_in_bits_cidx),
    .io__h2c_in_bits_port_id(tlb_io__h2c_in_bits_port_id),
    .io__h2c_in_bits_no_dma(tlb_io__h2c_in_bits_no_dma),
    .io__c2h_in_ready(tlb_io__c2h_in_ready),
    .io__c2h_in_valid(tlb_io__c2h_in_valid),
    .io__c2h_in_bits_addr(tlb_io__c2h_in_bits_addr),
    .io__c2h_in_bits_qid(tlb_io__c2h_in_bits_qid),
    .io__c2h_in_bits_error(tlb_io__c2h_in_bits_error),
    .io__c2h_in_bits_func(tlb_io__c2h_in_bits_func),
    .io__c2h_in_bits_port_id(tlb_io__c2h_in_bits_port_id),
    .io__c2h_in_bits_pfch_tag(tlb_io__c2h_in_bits_pfch_tag),
    .io__c2h_in_bits_len(tlb_io__c2h_in_bits_len),
    .io__h2c_out_ready(tlb_io__h2c_out_ready),
    .io__h2c_out_valid(tlb_io__h2c_out_valid),
    .io__h2c_out_bits_addr(tlb_io__h2c_out_bits_addr),
    .io__h2c_out_bits_len(tlb_io__h2c_out_bits_len),
    .io__h2c_out_bits_eop(tlb_io__h2c_out_bits_eop),
    .io__h2c_out_bits_sop(tlb_io__h2c_out_bits_sop),
    .io__h2c_out_bits_mrkr_req(tlb_io__h2c_out_bits_mrkr_req),
    .io__h2c_out_bits_sdi(tlb_io__h2c_out_bits_sdi),
    .io__h2c_out_bits_qid(tlb_io__h2c_out_bits_qid),
    .io__h2c_out_bits_error(tlb_io__h2c_out_bits_error),
    .io__h2c_out_bits_func(tlb_io__h2c_out_bits_func),
    .io__h2c_out_bits_cidx(tlb_io__h2c_out_bits_cidx),
    .io__h2c_out_bits_port_id(tlb_io__h2c_out_bits_port_id),
    .io__h2c_out_bits_no_dma(tlb_io__h2c_out_bits_no_dma),
    .io__c2h_out_ready(tlb_io__c2h_out_ready),
    .io__c2h_out_valid(tlb_io__c2h_out_valid),
    .io__c2h_out_bits_addr(tlb_io__c2h_out_bits_addr),
    .io__c2h_out_bits_qid(tlb_io__c2h_out_bits_qid),
    .io__c2h_out_bits_error(tlb_io__c2h_out_bits_error),
    .io__c2h_out_bits_func(tlb_io__c2h_out_bits_func),
    .io__c2h_out_bits_port_id(tlb_io__c2h_out_bits_port_id),
    .io__c2h_out_bits_pfch_tag(tlb_io__c2h_out_bits_pfch_tag),
    .io__c2h_out_bits_len(tlb_io__c2h_out_bits_len),
    .io__tlb_miss_count(tlb_io__tlb_miss_count),
    .io_tlb_miss_count(tlb_io_tlb_miss_count)
  );
  RegSlice_2 tlb_io_h2c_in_queue ( // @[RegSlices.scala 64:35]
    .clock(tlb_io_h2c_in_queue_clock),
    .reset(tlb_io_h2c_in_queue_reset),
    .io_upStream_ready(tlb_io_h2c_in_queue_io_upStream_ready),
    .io_upStream_valid(tlb_io_h2c_in_queue_io_upStream_valid),
    .io_upStream_bits_addr(tlb_io_h2c_in_queue_io_upStream_bits_addr),
    .io_upStream_bits_len(tlb_io_h2c_in_queue_io_upStream_bits_len),
    .io_upStream_bits_eop(tlb_io_h2c_in_queue_io_upStream_bits_eop),
    .io_upStream_bits_sop(tlb_io_h2c_in_queue_io_upStream_bits_sop),
    .io_upStream_bits_mrkr_req(tlb_io_h2c_in_queue_io_upStream_bits_mrkr_req),
    .io_upStream_bits_sdi(tlb_io_h2c_in_queue_io_upStream_bits_sdi),
    .io_upStream_bits_qid(tlb_io_h2c_in_queue_io_upStream_bits_qid),
    .io_upStream_bits_error(tlb_io_h2c_in_queue_io_upStream_bits_error),
    .io_upStream_bits_func(tlb_io_h2c_in_queue_io_upStream_bits_func),
    .io_upStream_bits_cidx(tlb_io_h2c_in_queue_io_upStream_bits_cidx),
    .io_upStream_bits_port_id(tlb_io_h2c_in_queue_io_upStream_bits_port_id),
    .io_upStream_bits_no_dma(tlb_io_h2c_in_queue_io_upStream_bits_no_dma),
    .io_downStream_ready(tlb_io_h2c_in_queue_io_downStream_ready),
    .io_downStream_valid(tlb_io_h2c_in_queue_io_downStream_valid),
    .io_downStream_bits_addr(tlb_io_h2c_in_queue_io_downStream_bits_addr),
    .io_downStream_bits_len(tlb_io_h2c_in_queue_io_downStream_bits_len),
    .io_downStream_bits_eop(tlb_io_h2c_in_queue_io_downStream_bits_eop),
    .io_downStream_bits_sop(tlb_io_h2c_in_queue_io_downStream_bits_sop),
    .io_downStream_bits_mrkr_req(tlb_io_h2c_in_queue_io_downStream_bits_mrkr_req),
    .io_downStream_bits_sdi(tlb_io_h2c_in_queue_io_downStream_bits_sdi),
    .io_downStream_bits_qid(tlb_io_h2c_in_queue_io_downStream_bits_qid),
    .io_downStream_bits_error(tlb_io_h2c_in_queue_io_downStream_bits_error),
    .io_downStream_bits_func(tlb_io_h2c_in_queue_io_downStream_bits_func),
    .io_downStream_bits_cidx(tlb_io_h2c_in_queue_io_downStream_bits_cidx),
    .io_downStream_bits_port_id(tlb_io_h2c_in_queue_io_downStream_bits_port_id),
    .io_downStream_bits_no_dma(tlb_io_h2c_in_queue_io_downStream_bits_no_dma)
  );
  RegSlice_3 tlb_io_c2h_in_queue ( // @[RegSlices.scala 64:35]
    .clock(tlb_io_c2h_in_queue_clock),
    .reset(tlb_io_c2h_in_queue_reset),
    .io_upStream_ready(tlb_io_c2h_in_queue_io_upStream_ready),
    .io_upStream_valid(tlb_io_c2h_in_queue_io_upStream_valid),
    .io_upStream_bits_addr(tlb_io_c2h_in_queue_io_upStream_bits_addr),
    .io_upStream_bits_qid(tlb_io_c2h_in_queue_io_upStream_bits_qid),
    .io_upStream_bits_error(tlb_io_c2h_in_queue_io_upStream_bits_error),
    .io_upStream_bits_func(tlb_io_c2h_in_queue_io_upStream_bits_func),
    .io_upStream_bits_port_id(tlb_io_c2h_in_queue_io_upStream_bits_port_id),
    .io_upStream_bits_pfch_tag(tlb_io_c2h_in_queue_io_upStream_bits_pfch_tag),
    .io_upStream_bits_len(tlb_io_c2h_in_queue_io_upStream_bits_len),
    .io_downStream_ready(tlb_io_c2h_in_queue_io_downStream_ready),
    .io_downStream_valid(tlb_io_c2h_in_queue_io_downStream_valid),
    .io_downStream_bits_addr(tlb_io_c2h_in_queue_io_downStream_bits_addr),
    .io_downStream_bits_qid(tlb_io_c2h_in_queue_io_downStream_bits_qid),
    .io_downStream_bits_error(tlb_io_c2h_in_queue_io_downStream_bits_error),
    .io_downStream_bits_func(tlb_io_c2h_in_queue_io_downStream_bits_func),
    .io_downStream_bits_port_id(tlb_io_c2h_in_queue_io_downStream_bits_port_id),
    .io_downStream_bits_pfch_tag(tlb_io_c2h_in_queue_io_downStream_bits_pfch_tag),
    .io_downStream_bits_len(tlb_io_c2h_in_queue_io_downStream_bits_len)
  );
  RegSlice_2 fifo_h2c_cmd_io_in_queue ( // @[RegSlices.scala 64:35]
    .clock(fifo_h2c_cmd_io_in_queue_clock),
    .reset(fifo_h2c_cmd_io_in_queue_reset),
    .io_upStream_ready(fifo_h2c_cmd_io_in_queue_io_upStream_ready),
    .io_upStream_valid(fifo_h2c_cmd_io_in_queue_io_upStream_valid),
    .io_upStream_bits_addr(fifo_h2c_cmd_io_in_queue_io_upStream_bits_addr),
    .io_upStream_bits_len(fifo_h2c_cmd_io_in_queue_io_upStream_bits_len),
    .io_upStream_bits_eop(fifo_h2c_cmd_io_in_queue_io_upStream_bits_eop),
    .io_upStream_bits_sop(fifo_h2c_cmd_io_in_queue_io_upStream_bits_sop),
    .io_upStream_bits_mrkr_req(fifo_h2c_cmd_io_in_queue_io_upStream_bits_mrkr_req),
    .io_upStream_bits_sdi(fifo_h2c_cmd_io_in_queue_io_upStream_bits_sdi),
    .io_upStream_bits_qid(fifo_h2c_cmd_io_in_queue_io_upStream_bits_qid),
    .io_upStream_bits_error(fifo_h2c_cmd_io_in_queue_io_upStream_bits_error),
    .io_upStream_bits_func(fifo_h2c_cmd_io_in_queue_io_upStream_bits_func),
    .io_upStream_bits_cidx(fifo_h2c_cmd_io_in_queue_io_upStream_bits_cidx),
    .io_upStream_bits_port_id(fifo_h2c_cmd_io_in_queue_io_upStream_bits_port_id),
    .io_upStream_bits_no_dma(fifo_h2c_cmd_io_in_queue_io_upStream_bits_no_dma),
    .io_downStream_ready(fifo_h2c_cmd_io_in_queue_io_downStream_ready),
    .io_downStream_valid(fifo_h2c_cmd_io_in_queue_io_downStream_valid),
    .io_downStream_bits_addr(fifo_h2c_cmd_io_in_queue_io_downStream_bits_addr),
    .io_downStream_bits_len(fifo_h2c_cmd_io_in_queue_io_downStream_bits_len),
    .io_downStream_bits_eop(fifo_h2c_cmd_io_in_queue_io_downStream_bits_eop),
    .io_downStream_bits_sop(fifo_h2c_cmd_io_in_queue_io_downStream_bits_sop),
    .io_downStream_bits_mrkr_req(fifo_h2c_cmd_io_in_queue_io_downStream_bits_mrkr_req),
    .io_downStream_bits_sdi(fifo_h2c_cmd_io_in_queue_io_downStream_bits_sdi),
    .io_downStream_bits_qid(fifo_h2c_cmd_io_in_queue_io_downStream_bits_qid),
    .io_downStream_bits_error(fifo_h2c_cmd_io_in_queue_io_downStream_bits_error),
    .io_downStream_bits_func(fifo_h2c_cmd_io_in_queue_io_downStream_bits_func),
    .io_downStream_bits_cidx(fifo_h2c_cmd_io_in_queue_io_downStream_bits_cidx),
    .io_downStream_bits_port_id(fifo_h2c_cmd_io_in_queue_io_downStream_bits_port_id),
    .io_downStream_bits_no_dma(fifo_h2c_cmd_io_in_queue_io_downStream_bits_no_dma)
  );
  PoorAXIL2Reg axil2reg ( // @[QDMADynamic.scala 86:76]
    .clock(axil2reg_clock),
    .reset(axil2reg_reset),
    .io_axi_aw_ready(axil2reg_io_axi_aw_ready),
    .io_axi_aw_valid(axil2reg_io_axi_aw_valid),
    .io_axi_aw_bits_addr(axil2reg_io_axi_aw_bits_addr),
    .io_axi_ar_ready(axil2reg_io_axi_ar_ready),
    .io_axi_ar_valid(axil2reg_io_axi_ar_valid),
    .io_axi_ar_bits_addr(axil2reg_io_axi_ar_bits_addr),
    .io_axi_w_ready(axil2reg_io_axi_w_ready),
    .io_axi_w_valid(axil2reg_io_axi_w_valid),
    .io_axi_w_bits_data(axil2reg_io_axi_w_bits_data),
    .io_axi_r_ready(axil2reg_io_axi_r_ready),
    .io_axi_r_valid(axil2reg_io_axi_r_valid),
    .io_axi_r_bits_data(axil2reg_io_axi_r_bits_data),
    .io_reg_control_0(axil2reg_io_reg_control_0),
    .io_reg_control_8(axil2reg_io_reg_control_8),
    .io_reg_control_9(axil2reg_io_reg_control_9),
    .io_reg_control_10(axil2reg_io_reg_control_10),
    .io_reg_control_11(axil2reg_io_reg_control_11),
    .io_reg_control_12(axil2reg_io_reg_control_12),
    .io_reg_control_13(axil2reg_io_reg_control_13),
    .io_reg_control_14(axil2reg_io_reg_control_14),
    .io_reg_status_300(axil2reg_io_reg_status_300),
    .io_reg_status_400(axil2reg_io_reg_status_400),
    .io_reg_status_401(axil2reg_io_reg_status_401),
    .io_reg_status_402(axil2reg_io_reg_status_402),
    .io_reg_status_403(axil2reg_io_reg_status_403),
    .io_reg_status_404(axil2reg_io_reg_status_404),
    .io_reg_status_405(axil2reg_io_reg_status_405),
    .io_reg_status_406(axil2reg_io_reg_status_406),
    .io_reg_status_407(axil2reg_io_reg_status_407),
    .io_reg_status_408(axil2reg_io_reg_status_408),
    .io_reg_status_409(axil2reg_io_reg_status_409),
    .io_reg_status_410(axil2reg_io_reg_status_410),
    .io_reg_status_411(axil2reg_io_reg_status_411),
    .io_reg_status_412(axil2reg_io_reg_status_412),
    .io_reg_status_413(axil2reg_io_reg_status_413),
    .io_reg_status_414(axil2reg_io_reg_status_414)
  );
  XConverter_4 io_axib_cvt_aw ( // @[XConverter.scala 61:33]
    .io_in_clk(io_axib_cvt_aw_io_in_clk),
    .io_out_clk(io_axib_cvt_aw_io_out_clk),
    .io_rstn(io_axib_cvt_aw_io_rstn),
    .io_in_ready(io_axib_cvt_aw_io_in_ready),
    .io_in_valid(io_axib_cvt_aw_io_in_valid),
    .io_in_bits_addr(io_axib_cvt_aw_io_in_bits_addr),
    .io_in_bits_burst(io_axib_cvt_aw_io_in_bits_burst),
    .io_in_bits_cache(io_axib_cvt_aw_io_in_bits_cache),
    .io_in_bits_id(io_axib_cvt_aw_io_in_bits_id),
    .io_in_bits_len(io_axib_cvt_aw_io_in_bits_len),
    .io_in_bits_lock(io_axib_cvt_aw_io_in_bits_lock),
    .io_in_bits_prot(io_axib_cvt_aw_io_in_bits_prot),
    .io_in_bits_size(io_axib_cvt_aw_io_in_bits_size),
    .io_out_ready(io_axib_cvt_aw_io_out_ready),
    .io_out_valid(io_axib_cvt_aw_io_out_valid),
    .io_out_bits_addr(io_axib_cvt_aw_io_out_bits_addr)
  );
  XConverter_4 io_axib_cvt_ar ( // @[XConverter.scala 61:33]
    .io_in_clk(io_axib_cvt_ar_io_in_clk),
    .io_out_clk(io_axib_cvt_ar_io_out_clk),
    .io_rstn(io_axib_cvt_ar_io_rstn),
    .io_in_ready(io_axib_cvt_ar_io_in_ready),
    .io_in_valid(io_axib_cvt_ar_io_in_valid),
    .io_in_bits_addr(io_axib_cvt_ar_io_in_bits_addr),
    .io_in_bits_burst(io_axib_cvt_ar_io_in_bits_burst),
    .io_in_bits_cache(io_axib_cvt_ar_io_in_bits_cache),
    .io_in_bits_id(io_axib_cvt_ar_io_in_bits_id),
    .io_in_bits_len(io_axib_cvt_ar_io_in_bits_len),
    .io_in_bits_lock(io_axib_cvt_ar_io_in_bits_lock),
    .io_in_bits_prot(io_axib_cvt_ar_io_in_bits_prot),
    .io_in_bits_size(io_axib_cvt_ar_io_in_bits_size),
    .io_out_ready(io_axib_cvt_ar_io_out_ready),
    .io_out_valid(io_axib_cvt_ar_io_out_valid),
    .io_out_bits_addr(io_axib_cvt_ar_io_out_bits_addr)
  );
  XConverter_6 io_axib_cvt_w ( // @[XConverter.scala 61:33]
    .io_in_clk(io_axib_cvt_w_io_in_clk),
    .io_out_clk(io_axib_cvt_w_io_out_clk),
    .io_rstn(io_axib_cvt_w_io_rstn),
    .io_in_ready(io_axib_cvt_w_io_in_ready),
    .io_in_valid(io_axib_cvt_w_io_in_valid),
    .io_in_bits_data(io_axib_cvt_w_io_in_bits_data),
    .io_in_bits_last(io_axib_cvt_w_io_in_bits_last),
    .io_in_bits_strb(io_axib_cvt_w_io_in_bits_strb),
    .io_out_ready(io_axib_cvt_w_io_out_ready),
    .io_out_valid(io_axib_cvt_w_io_out_valid),
    .io_out_bits_data(io_axib_cvt_w_io_out_bits_data)
  );
  XConverter_7 io_axib_cvt_r ( // @[XConverter.scala 61:33]
    .io_in_clk(io_axib_cvt_r_io_in_clk),
    .io_out_clk(io_axib_cvt_r_io_out_clk),
    .io_rstn(io_axib_cvt_r_io_rstn),
    .io_in_ready(io_axib_cvt_r_io_in_ready),
    .io_in_bits_data(io_axib_cvt_r_io_in_bits_data),
    .io_out_ready(io_axib_cvt_r_io_out_ready),
    .io_out_valid(io_axib_cvt_r_io_out_valid),
    .io_out_bits_data(io_axib_cvt_r_io_out_bits_data),
    .io_out_bits_last(io_axib_cvt_r_io_out_bits_last),
    .io_out_bits_resp(io_axib_cvt_r_io_out_bits_resp),
    .io_out_bits_id(io_axib_cvt_r_io_out_bits_id)
  );
  XConverter_8 io_axib_cvt_b ( // @[XConverter.scala 61:33]
    .io_in_clk(io_axib_cvt_b_io_in_clk),
    .io_out_clk(io_axib_cvt_b_io_out_clk),
    .io_rstn(io_axib_cvt_b_io_rstn),
    .io_out_ready(io_axib_cvt_b_io_out_ready),
    .io_out_valid(io_axib_cvt_b_io_out_valid),
    .io_out_bits_id(io_axib_cvt_b_io_out_bits_id),
    .io_out_bits_resp(io_axib_cvt_b_io_out_bits_resp)
  );
  XConverter_9 axil2reg_io_axi_cvt_aw ( // @[XConverter.scala 61:33]
    .io_in_clk(axil2reg_io_axi_cvt_aw_io_in_clk),
    .io_out_clk(axil2reg_io_axi_cvt_aw_io_out_clk),
    .io_rstn(axil2reg_io_axi_cvt_aw_io_rstn),
    .io_in_ready(axil2reg_io_axi_cvt_aw_io_in_ready),
    .io_in_valid(axil2reg_io_axi_cvt_aw_io_in_valid),
    .io_in_bits_addr(axil2reg_io_axi_cvt_aw_io_in_bits_addr),
    .io_out_ready(axil2reg_io_axi_cvt_aw_io_out_ready),
    .io_out_valid(axil2reg_io_axi_cvt_aw_io_out_valid),
    .io_out_bits_addr(axil2reg_io_axi_cvt_aw_io_out_bits_addr)
  );
  XConverter_9 axil2reg_io_axi_cvt_ar ( // @[XConverter.scala 61:33]
    .io_in_clk(axil2reg_io_axi_cvt_ar_io_in_clk),
    .io_out_clk(axil2reg_io_axi_cvt_ar_io_out_clk),
    .io_rstn(axil2reg_io_axi_cvt_ar_io_rstn),
    .io_in_ready(axil2reg_io_axi_cvt_ar_io_in_ready),
    .io_in_valid(axil2reg_io_axi_cvt_ar_io_in_valid),
    .io_in_bits_addr(axil2reg_io_axi_cvt_ar_io_in_bits_addr),
    .io_out_ready(axil2reg_io_axi_cvt_ar_io_out_ready),
    .io_out_valid(axil2reg_io_axi_cvt_ar_io_out_valid),
    .io_out_bits_addr(axil2reg_io_axi_cvt_ar_io_out_bits_addr)
  );
  XConverter_11 axil2reg_io_axi_cvt_w ( // @[XConverter.scala 61:33]
    .io_in_clk(axil2reg_io_axi_cvt_w_io_in_clk),
    .io_out_clk(axil2reg_io_axi_cvt_w_io_out_clk),
    .io_rstn(axil2reg_io_axi_cvt_w_io_rstn),
    .io_in_ready(axil2reg_io_axi_cvt_w_io_in_ready),
    .io_in_valid(axil2reg_io_axi_cvt_w_io_in_valid),
    .io_in_bits_data(axil2reg_io_axi_cvt_w_io_in_bits_data),
    .io_in_bits_strb(axil2reg_io_axi_cvt_w_io_in_bits_strb),
    .io_out_ready(axil2reg_io_axi_cvt_w_io_out_ready),
    .io_out_valid(axil2reg_io_axi_cvt_w_io_out_valid),
    .io_out_bits_data(axil2reg_io_axi_cvt_w_io_out_bits_data)
  );
  XConverter_12 axil2reg_io_axi_cvt_r ( // @[XConverter.scala 61:33]
    .io_in_clk(axil2reg_io_axi_cvt_r_io_in_clk),
    .io_out_clk(axil2reg_io_axi_cvt_r_io_out_clk),
    .io_rstn(axil2reg_io_axi_cvt_r_io_rstn),
    .io_in_ready(axil2reg_io_axi_cvt_r_io_in_ready),
    .io_in_valid(axil2reg_io_axi_cvt_r_io_in_valid),
    .io_in_bits_data(axil2reg_io_axi_cvt_r_io_in_bits_data),
    .io_out_ready(axil2reg_io_axi_cvt_r_io_out_ready),
    .io_out_valid(axil2reg_io_axi_cvt_r_io_out_valid),
    .io_out_bits_data(axil2reg_io_axi_cvt_r_io_out_bits_data),
    .io_out_bits_resp(axil2reg_io_axi_cvt_r_io_out_bits_resp)
  );
  XConverter_13 axil2reg_io_axi_cvt_b ( // @[XConverter.scala 61:33]
    .io_in_clk(axil2reg_io_axi_cvt_b_io_in_clk),
    .io_out_clk(axil2reg_io_axi_cvt_b_io_out_clk),
    .io_rstn(axil2reg_io_axi_cvt_b_io_rstn),
    .io_out_ready(axil2reg_io_axi_cvt_b_io_out_ready),
    .io_out_valid(axil2reg_io_axi_cvt_b_io_out_valid),
    .io_out_bits_resp(axil2reg_io_axi_cvt_b_io_out_bits_resp)
  );
  DataBoundarySplit boundary_split ( // @[QDMADynamic.scala 116:82]
    .clock(boundary_split_clock),
    .reset(boundary_split_reset),
    .io_cmd_in_ready(boundary_split_io_cmd_in_ready),
    .io_cmd_in_valid(boundary_split_io_cmd_in_valid),
    .io_cmd_in_bits_addr(boundary_split_io_cmd_in_bits_addr),
    .io_cmd_in_bits_qid(boundary_split_io_cmd_in_bits_qid),
    .io_cmd_in_bits_error(boundary_split_io_cmd_in_bits_error),
    .io_cmd_in_bits_func(boundary_split_io_cmd_in_bits_func),
    .io_cmd_in_bits_port_id(boundary_split_io_cmd_in_bits_port_id),
    .io_cmd_in_bits_pfch_tag(boundary_split_io_cmd_in_bits_pfch_tag),
    .io_cmd_in_bits_len(boundary_split_io_cmd_in_bits_len),
    .io_data_out_ready(boundary_split_io_data_out_ready),
    .io_data_out_valid(boundary_split_io_data_out_valid),
    .io_data_out_bits_data(boundary_split_io_data_out_bits_data),
    .io_data_out_bits_tcrc(boundary_split_io_data_out_bits_tcrc),
    .io_data_out_bits_ctrl_marker(boundary_split_io_data_out_bits_ctrl_marker),
    .io_data_out_bits_ctrl_ecc(boundary_split_io_data_out_bits_ctrl_ecc),
    .io_data_out_bits_ctrl_len(boundary_split_io_data_out_bits_ctrl_len),
    .io_data_out_bits_ctrl_port_id(boundary_split_io_data_out_bits_ctrl_port_id),
    .io_data_out_bits_ctrl_qid(boundary_split_io_data_out_bits_ctrl_qid),
    .io_data_out_bits_ctrl_has_cmpt(boundary_split_io_data_out_bits_ctrl_has_cmpt),
    .io_data_out_bits_last(boundary_split_io_data_out_bits_last),
    .io_data_out_bits_mty(boundary_split_io_data_out_bits_mty),
    .io_cmd_out_ready(boundary_split_io_cmd_out_ready),
    .io_cmd_out_valid(boundary_split_io_cmd_out_valid),
    .io_cmd_out_bits_addr(boundary_split_io_cmd_out_bits_addr),
    .io_cmd_out_bits_qid(boundary_split_io_cmd_out_bits_qid),
    .io_cmd_out_bits_error(boundary_split_io_cmd_out_bits_error),
    .io_cmd_out_bits_func(boundary_split_io_cmd_out_bits_func),
    .io_cmd_out_bits_port_id(boundary_split_io_cmd_out_bits_port_id),
    .io_cmd_out_bits_pfch_tag(boundary_split_io_cmd_out_bits_pfch_tag),
    .io_cmd_out_bits_len(boundary_split_io_cmd_out_bits_len)
  );
  assign io_qdma_port_m_axib_awready = io_axib_cvt_aw_io_in_ready; // @[QDMADynamic.scala 92:24 XConverter.scala 35:33]
  assign io_qdma_port_m_axib_wready = io_axib_cvt_w_io_in_ready; // @[QDMADynamic.scala 92:24 XConverter.scala 37:33]
  assign io_qdma_port_m_axib_bid = io_axib_cvt_b_io_out_bits_id; // @[QDMADynamic.scala 92:24 XConverter.scala 39:33]
  assign io_qdma_port_m_axib_bresp = io_axib_cvt_b_io_out_bits_resp; // @[QDMADynamic.scala 92:24 XConverter.scala 39:33]
  assign io_qdma_port_m_axib_bvalid = io_axib_cvt_b_io_out_valid; // @[QDMADynamic.scala 92:24 XConverter.scala 39:33]
  assign io_qdma_port_m_axib_arready = io_axib_cvt_ar_io_in_ready; // @[QDMADynamic.scala 92:24 XConverter.scala 36:33]
  assign io_qdma_port_m_axib_rid = io_axib_cvt_r_io_out_bits_id; // @[QDMADynamic.scala 92:24 XConverter.scala 38:33]
  assign io_qdma_port_m_axib_rdata = io_axib_cvt_r_io_out_bits_data; // @[QDMADynamic.scala 92:24 XConverter.scala 38:33]
  assign io_qdma_port_m_axib_rresp = io_axib_cvt_r_io_out_bits_resp; // @[QDMADynamic.scala 92:24 XConverter.scala 38:33]
  assign io_qdma_port_m_axib_rlast = io_axib_cvt_r_io_out_bits_last; // @[QDMADynamic.scala 92:24 XConverter.scala 38:33]
  assign io_qdma_port_m_axib_rvalid = io_axib_cvt_r_io_out_valid; // @[QDMADynamic.scala 92:24 XConverter.scala 38:33]
  assign io_qdma_port_m_axil_awready = axil2reg_io_axi_cvt_aw_io_in_ready; // @[QDMADynamic.scala 107:24 XConverter.scala 35:33]
  assign io_qdma_port_m_axil_wready = axil2reg_io_axi_cvt_w_io_in_ready; // @[QDMADynamic.scala 107:24 XConverter.scala 37:33]
  assign io_qdma_port_m_axil_bresp = axil2reg_io_axi_cvt_b_io_out_bits_resp; // @[QDMADynamic.scala 107:24 XConverter.scala 39:33]
  assign io_qdma_port_m_axil_bvalid = axil2reg_io_axi_cvt_b_io_out_valid; // @[QDMADynamic.scala 107:24 XConverter.scala 39:33]
  assign io_qdma_port_m_axil_arready = axil2reg_io_axi_cvt_ar_io_in_ready; // @[QDMADynamic.scala 107:24 XConverter.scala 36:33]
  assign io_qdma_port_m_axil_rdata = axil2reg_io_axi_cvt_r_io_out_bits_data; // @[QDMADynamic.scala 107:24 XConverter.scala 38:33]
  assign io_qdma_port_m_axil_rresp = axil2reg_io_axi_cvt_r_io_out_bits_resp; // @[QDMADynamic.scala 107:24 XConverter.scala 38:33]
  assign io_qdma_port_m_axil_rvalid = axil2reg_io_axi_cvt_r_io_out_valid; // @[QDMADynamic.scala 107:24 XConverter.scala 38:33]
  assign io_qdma_port_h2c_byp_in_st_addr = fifo_h2c_cmd_out_queue_io_downStream_bits_addr; // @[RegSlices.scala 63:38 RegSlices.scala 66:41]
  assign io_qdma_port_h2c_byp_in_st_len = fifo_h2c_cmd_out_queue_io_downStream_bits_len; // @[RegSlices.scala 63:38 RegSlices.scala 66:41]
  assign io_qdma_port_h2c_byp_in_st_eop = fifo_h2c_cmd_out_queue_io_downStream_bits_eop; // @[RegSlices.scala 63:38 RegSlices.scala 66:41]
  assign io_qdma_port_h2c_byp_in_st_sop = fifo_h2c_cmd_out_queue_io_downStream_bits_sop; // @[RegSlices.scala 63:38 RegSlices.scala 66:41]
  assign io_qdma_port_h2c_byp_in_st_mrkr_req = fifo_h2c_cmd_out_queue_io_downStream_bits_mrkr_req; // @[RegSlices.scala 63:38 RegSlices.scala 66:41]
  assign io_qdma_port_h2c_byp_in_st_sdi = fifo_h2c_cmd_out_queue_io_downStream_bits_sdi; // @[RegSlices.scala 63:38 RegSlices.scala 66:41]
  assign io_qdma_port_h2c_byp_in_st_qid = fifo_h2c_cmd_out_queue_io_downStream_bits_qid; // @[RegSlices.scala 63:38 RegSlices.scala 66:41]
  assign io_qdma_port_h2c_byp_in_st_error = fifo_h2c_cmd_out_queue_io_downStream_bits_error; // @[RegSlices.scala 63:38 RegSlices.scala 66:41]
  assign io_qdma_port_h2c_byp_in_st_func = fifo_h2c_cmd_out_queue_io_downStream_bits_func; // @[RegSlices.scala 63:38 RegSlices.scala 66:41]
  assign io_qdma_port_h2c_byp_in_st_cidx = fifo_h2c_cmd_out_queue_io_downStream_bits_cidx; // @[RegSlices.scala 63:38 RegSlices.scala 66:41]
  assign io_qdma_port_h2c_byp_in_st_port_id = fifo_h2c_cmd_out_queue_io_downStream_bits_port_id; // @[RegSlices.scala 63:38 RegSlices.scala 66:41]
  assign io_qdma_port_h2c_byp_in_st_no_dma = fifo_h2c_cmd_out_queue_io_downStream_bits_no_dma; // @[RegSlices.scala 63:38 RegSlices.scala 66:41]
  assign io_qdma_port_h2c_byp_in_st_vld = fifo_h2c_cmd_out_queue_io_downStream_valid; // @[RegSlices.scala 63:38 RegSlices.scala 66:41]
  assign io_qdma_port_c2h_byp_in_st_csh_addr = fifo_c2h_cmd_out_queue_io_downStream_bits_addr; // @[RegSlices.scala 63:38 RegSlices.scala 66:41]
  assign io_qdma_port_c2h_byp_in_st_csh_qid = fifo_c2h_cmd_out_queue_io_downStream_bits_qid; // @[RegSlices.scala 63:38 RegSlices.scala 66:41]
  assign io_qdma_port_c2h_byp_in_st_csh_error = fifo_c2h_cmd_out_queue_io_downStream_bits_error; // @[RegSlices.scala 63:38 RegSlices.scala 66:41]
  assign io_qdma_port_c2h_byp_in_st_csh_func = fifo_c2h_cmd_out_queue_io_downStream_bits_func; // @[RegSlices.scala 63:38 RegSlices.scala 66:41]
  assign io_qdma_port_c2h_byp_in_st_csh_port_id = fifo_c2h_cmd_out_queue_io_downStream_bits_port_id; // @[RegSlices.scala 63:38 RegSlices.scala 66:41]
  assign io_qdma_port_c2h_byp_in_st_csh_pfch_tag = fifo_c2h_cmd_out_queue_io_downStream_bits_pfch_tag; // @[RegSlices.scala 63:38 RegSlices.scala 66:41]
  assign io_qdma_port_c2h_byp_in_st_csh_vld = fifo_c2h_cmd_out_queue_io_downStream_valid; // @[RegSlices.scala 63:38 RegSlices.scala 66:41]
  assign io_qdma_port_s_axis_c2h_tdata = fifo_c2h_data_out_queue_io_downStream_bits_data; // @[RegSlices.scala 63:38 RegSlices.scala 66:41]
  assign io_qdma_port_s_axis_c2h_tcrc = fifo_c2h_data_out_queue_io_downStream_bits_tcrc; // @[RegSlices.scala 63:38 RegSlices.scala 66:41]
  assign io_qdma_port_s_axis_c2h_ctrl_marker = fifo_c2h_data_out_queue_io_downStream_bits_ctrl_marker; // @[RegSlices.scala 63:38 RegSlices.scala 66:41]
  assign io_qdma_port_s_axis_c2h_ctrl_ecc = fifo_c2h_data_out_queue_io_downStream_bits_ctrl_ecc; // @[RegSlices.scala 63:38 RegSlices.scala 66:41]
  assign io_qdma_port_s_axis_c2h_ctrl_len = fifo_c2h_data_out_queue_io_downStream_bits_ctrl_len; // @[RegSlices.scala 63:38 RegSlices.scala 66:41]
  assign io_qdma_port_s_axis_c2h_ctrl_port_id = fifo_c2h_data_out_queue_io_downStream_bits_ctrl_port_id; // @[RegSlices.scala 63:38 RegSlices.scala 66:41]
  assign io_qdma_port_s_axis_c2h_ctrl_qid = fifo_c2h_data_out_queue_io_downStream_bits_ctrl_qid; // @[RegSlices.scala 63:38 RegSlices.scala 66:41]
  assign io_qdma_port_s_axis_c2h_ctrl_has_cmpt = fifo_c2h_data_out_queue_io_downStream_bits_ctrl_has_cmpt; // @[RegSlices.scala 63:38 RegSlices.scala 66:41]
  assign io_qdma_port_s_axis_c2h_mty = fifo_c2h_data_out_queue_io_downStream_bits_mty; // @[RegSlices.scala 63:38 RegSlices.scala 66:41]
  assign io_qdma_port_s_axis_c2h_tlast = fifo_c2h_data_out_queue_io_downStream_bits_last; // @[RegSlices.scala 63:38 RegSlices.scala 66:41]
  assign io_qdma_port_s_axis_c2h_tvalid = fifo_c2h_data_out_queue_io_downStream_valid; // @[RegSlices.scala 63:38 RegSlices.scala 66:41]
  assign io_qdma_port_m_axis_h2c_tready = fifo_h2c_data_io_in_queue_io_upStream_ready; // @[QDMADynamic.scala 50:39 RegSlices.scala 65:41]
  assign io_h2c_cmd_ready = check_h2c_io_in_queue_io_upStream_ready; // @[RegSlices.scala 65:41]
  assign io_h2c_data_valid = fifo_h2c_data_io__out_valid; // @[QDMADynamic.scala 53:33]
  assign io_reg_control_0 = axil2reg_io_reg_control_0; // @[QDMADynamic.scala 89:33]
  assign io_reg_control_8 = axil2reg_io_reg_control_8; // @[QDMADynamic.scala 89:33]
  assign io_reg_control_9 = axil2reg_io_reg_control_9; // @[QDMADynamic.scala 89:33]
  assign io_reg_control_10 = axil2reg_io_reg_control_10; // @[QDMADynamic.scala 89:33]
  assign io_reg_control_11 = axil2reg_io_reg_control_11; // @[QDMADynamic.scala 89:33]
  assign io_reg_control_12 = axil2reg_io_reg_control_12; // @[QDMADynamic.scala 89:33]
  assign io_reg_control_13 = axil2reg_io_reg_control_13; // @[QDMADynamic.scala 89:33]
  assign io_reg_control_14 = axil2reg_io_reg_control_14; // @[QDMADynamic.scala 89:33]
  assign io_axib_aw_valid = io_axib_cvt_aw_io_out_valid; // @[XConverter.scala 22:39 XConverter.scala 41:33]
  assign io_axib_aw_bits_addr = io_axib_cvt_aw_io_out_bits_addr; // @[XConverter.scala 22:39 XConverter.scala 41:33]
  assign io_axib_w_valid = io_axib_cvt_w_io_out_valid; // @[XConverter.scala 22:39 XConverter.scala 43:33]
  assign io_axib_w_bits_data = io_axib_cvt_w_io_out_bits_data; // @[XConverter.scala 22:39 XConverter.scala 43:33]
  assign io_axib_r_ready = io_axib_cvt_r_io_in_ready; // @[XConverter.scala 22:39 XConverter.scala 44:41]
  assign io_out_valid = fifo_h2c_cmd_io_out_valid;
  assign counter_4_0 = counter_4;
  assign io_out_ready = fifo_c2h_data_io_out_ready;
  assign counter_7_0 = counter_7;
  assign counter_1_0 = counter_1;
  assign io_in_ready = fifo_h2c_data_io_in_ready;
  assign counter_3_1 = counter_3;
  assign io_out_ready_0 = fifo_c2h_cmd_io_out_ready_0;
  assign counter_6_0 = counter_6;
  assign io_out_valid_0 = fifo_c2h_data_io_out_valid_0;
  assign counter_0 = counter;
  assign io_in_valid = fifo_h2c_data_io_in_valid;
  assign io_tlb_miss_count = tlb_io_tlb_miss_count;
  assign io_out_valid_1 = fifo_c2h_cmd_io_out_valid_1;
  assign counter_2_1 = counter_2;
  assign counter_5_0 = counter_5;
  assign io_out_ready_1 = fifo_h2c_cmd_io_out_ready_1;
  assign sw_reset_pad_I = io_reg_control_14[0]; // @[QDMADynamic.scala 45:51]
  assign fifo_h2c_data_io__in_clk = io_qdma_port_axi_aclk; // @[QDMADynamic.scala 47:53]
  assign fifo_h2c_data_io__out_clk = io_user_clk; // @[XConverter.scala 63:33]
  assign fifo_h2c_data_io__rstn = io_qdma_port_axi_aresetn; // @[QDMADynamic.scala 48:51]
  assign fifo_h2c_data_io__in_valid = fifo_h2c_data_io_in_queue_io_downStream_valid; // @[RegSlices.scala 63:38 RegSlices.scala 66:41]
  assign fifo_h2c_data_io__in_bits_data = fifo_h2c_data_io_in_queue_io_downStream_bits_data; // @[RegSlices.scala 63:38 RegSlices.scala 66:41]
  assign fifo_h2c_data_io__in_bits_tcrc = fifo_h2c_data_io_in_queue_io_downStream_bits_tcrc; // @[RegSlices.scala 63:38 RegSlices.scala 66:41]
  assign fifo_h2c_data_io__in_bits_tuser_qid = fifo_h2c_data_io_in_queue_io_downStream_bits_tuser_qid; // @[RegSlices.scala 63:38 RegSlices.scala 66:41]
  assign fifo_h2c_data_io__in_bits_tuser_port_id = fifo_h2c_data_io_in_queue_io_downStream_bits_tuser_port_id; // @[RegSlices.scala 63:38 RegSlices.scala 66:41]
  assign fifo_h2c_data_io__in_bits_tuser_err = fifo_h2c_data_io_in_queue_io_downStream_bits_tuser_err; // @[RegSlices.scala 63:38 RegSlices.scala 66:41]
  assign fifo_h2c_data_io__in_bits_tuser_mdata = fifo_h2c_data_io_in_queue_io_downStream_bits_tuser_mdata; // @[RegSlices.scala 63:38 RegSlices.scala 66:41]
  assign fifo_h2c_data_io__in_bits_tuser_mty = fifo_h2c_data_io_in_queue_io_downStream_bits_tuser_mty; // @[RegSlices.scala 63:38 RegSlices.scala 66:41]
  assign fifo_h2c_data_io__in_bits_tuser_zero_byte = fifo_h2c_data_io_in_queue_io_downStream_bits_tuser_zero_byte; // @[RegSlices.scala 63:38 RegSlices.scala 66:41]
  assign fifo_h2c_data_io__in_bits_last = fifo_h2c_data_io_in_queue_io_downStream_bits_last; // @[RegSlices.scala 63:38 RegSlices.scala 66:41]
  assign fifo_h2c_data_io_in_queue_clock = io_qdma_port_axi_aclk; // @[QDMADynamic.scala 47:53]
  assign fifo_h2c_data_io_in_queue_reset = ~io_qdma_port_axi_aresetn; // @[QDMADynamic.scala 52:73]
  assign fifo_h2c_data_io_in_queue_io_upStream_valid = io_qdma_port_m_axis_h2c_tvalid; // @[QDMADynamic.scala 50:39 QDMADynamic.scala 201:57]
  assign fifo_h2c_data_io_in_queue_io_upStream_bits_data = io_qdma_port_m_axis_h2c_tdata; // @[QDMADynamic.scala 50:39 QDMADynamic.scala 192:57]
  assign fifo_h2c_data_io_in_queue_io_upStream_bits_tcrc = io_qdma_port_m_axis_h2c_tcrc; // @[QDMADynamic.scala 50:39 QDMADynamic.scala 193:57]
  assign fifo_h2c_data_io_in_queue_io_upStream_bits_tuser_qid = io_qdma_port_m_axis_h2c_tuser_qid; // @[QDMADynamic.scala 50:39 QDMADynamic.scala 194:57]
  assign fifo_h2c_data_io_in_queue_io_upStream_bits_tuser_port_id = io_qdma_port_m_axis_h2c_tuser_port_id; // @[QDMADynamic.scala 50:39 QDMADynamic.scala 195:49]
  assign fifo_h2c_data_io_in_queue_io_upStream_bits_tuser_err = io_qdma_port_m_axis_h2c_tuser_err; // @[QDMADynamic.scala 50:39 QDMADynamic.scala 196:57]
  assign fifo_h2c_data_io_in_queue_io_upStream_bits_tuser_mdata = io_qdma_port_m_axis_h2c_tuser_mdata; // @[QDMADynamic.scala 50:39 QDMADynamic.scala 197:57]
  assign fifo_h2c_data_io_in_queue_io_upStream_bits_tuser_mty = io_qdma_port_m_axis_h2c_tuser_mty; // @[QDMADynamic.scala 50:39 QDMADynamic.scala 198:57]
  assign fifo_h2c_data_io_in_queue_io_upStream_bits_tuser_zero_byte = io_qdma_port_m_axis_h2c_tuser_zero_byte; // @[QDMADynamic.scala 50:39 QDMADynamic.scala 199:49]
  assign fifo_h2c_data_io_in_queue_io_upStream_bits_last = io_qdma_port_m_axis_h2c_tlast; // @[QDMADynamic.scala 50:39 QDMADynamic.scala 200:57]
  assign fifo_h2c_data_io_in_queue_io_downStream_ready = fifo_h2c_data_io__in_ready; // @[RegSlices.scala 63:38 QDMADynamic.scala 52:41]
  assign fifo_c2h_data_io__in_clk = io_user_clk; // @[XConverter.scala 62:33]
  assign fifo_c2h_data_io__out_clk = io_qdma_port_axi_aclk; // @[QDMADynamic.scala 47:53]
  assign fifo_c2h_data_io__rstn = io_user_arstn; // @[XConverter.scala 64:41]
  assign fifo_c2h_data_io__in_valid = boundary_split_io_data_out_valid; // @[QDMADynamic.scala 120:41]
  assign fifo_c2h_data_io__in_bits_data = boundary_split_io_data_out_bits_data; // @[QDMADynamic.scala 120:41]
  assign fifo_c2h_data_io__in_bits_tcrc = boundary_split_io_data_out_bits_tcrc; // @[QDMADynamic.scala 120:41]
  assign fifo_c2h_data_io__in_bits_ctrl_marker = boundary_split_io_data_out_bits_ctrl_marker; // @[QDMADynamic.scala 120:41]
  assign fifo_c2h_data_io__in_bits_ctrl_ecc = boundary_split_io_data_out_bits_ctrl_ecc; // @[QDMADynamic.scala 120:41]
  assign fifo_c2h_data_io__in_bits_ctrl_len = boundary_split_io_data_out_bits_ctrl_len; // @[QDMADynamic.scala 120:41]
  assign fifo_c2h_data_io__in_bits_ctrl_port_id = boundary_split_io_data_out_bits_ctrl_port_id; // @[QDMADynamic.scala 120:41]
  assign fifo_c2h_data_io__in_bits_ctrl_qid = boundary_split_io_data_out_bits_ctrl_qid; // @[QDMADynamic.scala 120:41]
  assign fifo_c2h_data_io__in_bits_ctrl_has_cmpt = boundary_split_io_data_out_bits_ctrl_has_cmpt; // @[QDMADynamic.scala 120:41]
  assign fifo_c2h_data_io__in_bits_last = boundary_split_io_data_out_bits_last; // @[QDMADynamic.scala 120:41]
  assign fifo_c2h_data_io__in_bits_mty = boundary_split_io_data_out_bits_mty; // @[QDMADynamic.scala 120:41]
  assign fifo_c2h_data_io__out_ready = fifo_c2h_data_out_queue_io_upStream_ready; // @[RegSlices.scala 65:41]
  assign fifo_c2h_data_out_queue_clock = io_qdma_port_axi_aclk; // @[QDMADynamic.scala 47:53]
  assign fifo_c2h_data_out_queue_reset = ~io_qdma_port_axi_aresetn; // @[QDMADynamic.scala 56:64]
  assign fifo_c2h_data_out_queue_io_upStream_valid = fifo_c2h_data_io__out_valid; // @[RegSlices.scala 65:41]
  assign fifo_c2h_data_out_queue_io_upStream_bits_data = fifo_c2h_data_io__out_bits_data; // @[RegSlices.scala 65:41]
  assign fifo_c2h_data_out_queue_io_upStream_bits_tcrc = fifo_c2h_data_io__out_bits_tcrc; // @[RegSlices.scala 65:41]
  assign fifo_c2h_data_out_queue_io_upStream_bits_ctrl_marker = fifo_c2h_data_io__out_bits_ctrl_marker; // @[RegSlices.scala 65:41]
  assign fifo_c2h_data_out_queue_io_upStream_bits_ctrl_ecc = fifo_c2h_data_io__out_bits_ctrl_ecc; // @[RegSlices.scala 65:41]
  assign fifo_c2h_data_out_queue_io_upStream_bits_ctrl_len = fifo_c2h_data_io__out_bits_ctrl_len; // @[RegSlices.scala 65:41]
  assign fifo_c2h_data_out_queue_io_upStream_bits_ctrl_port_id = fifo_c2h_data_io__out_bits_ctrl_port_id; // @[RegSlices.scala 65:41]
  assign fifo_c2h_data_out_queue_io_upStream_bits_ctrl_qid = fifo_c2h_data_io__out_bits_ctrl_qid; // @[RegSlices.scala 65:41]
  assign fifo_c2h_data_out_queue_io_upStream_bits_ctrl_has_cmpt = fifo_c2h_data_io__out_bits_ctrl_has_cmpt; // @[RegSlices.scala 65:41]
  assign fifo_c2h_data_out_queue_io_upStream_bits_last = fifo_c2h_data_io__out_bits_last; // @[RegSlices.scala 65:41]
  assign fifo_c2h_data_out_queue_io_upStream_bits_mty = fifo_c2h_data_io__out_bits_mty; // @[RegSlices.scala 65:41]
  assign fifo_c2h_data_out_queue_io_downStream_ready = io_qdma_port_s_axis_c2h_tready; // @[RegSlices.scala 63:38 QDMADynamic.scala 189:57]
  assign fifo_h2c_cmd_io__in_clk = io_user_clk; // @[XConverter.scala 62:33]
  assign fifo_h2c_cmd_io__out_clk = io_qdma_port_axi_aclk; // @[QDMADynamic.scala 47:53]
  assign fifo_h2c_cmd_io__rstn = io_user_arstn; // @[XConverter.scala 64:41]
  assign fifo_h2c_cmd_io__in_valid = fifo_h2c_cmd_io_in_queue_io_downStream_valid; // @[RegSlices.scala 63:38 RegSlices.scala 66:41]
  assign fifo_h2c_cmd_io__in_bits_addr = fifo_h2c_cmd_io_in_queue_io_downStream_bits_addr; // @[RegSlices.scala 63:38 RegSlices.scala 66:41]
  assign fifo_h2c_cmd_io__in_bits_len = fifo_h2c_cmd_io_in_queue_io_downStream_bits_len; // @[RegSlices.scala 63:38 RegSlices.scala 66:41]
  assign fifo_h2c_cmd_io__in_bits_eop = fifo_h2c_cmd_io_in_queue_io_downStream_bits_eop; // @[RegSlices.scala 63:38 RegSlices.scala 66:41]
  assign fifo_h2c_cmd_io__in_bits_sop = fifo_h2c_cmd_io_in_queue_io_downStream_bits_sop; // @[RegSlices.scala 63:38 RegSlices.scala 66:41]
  assign fifo_h2c_cmd_io__in_bits_mrkr_req = fifo_h2c_cmd_io_in_queue_io_downStream_bits_mrkr_req; // @[RegSlices.scala 63:38 RegSlices.scala 66:41]
  assign fifo_h2c_cmd_io__in_bits_sdi = fifo_h2c_cmd_io_in_queue_io_downStream_bits_sdi; // @[RegSlices.scala 63:38 RegSlices.scala 66:41]
  assign fifo_h2c_cmd_io__in_bits_qid = fifo_h2c_cmd_io_in_queue_io_downStream_bits_qid; // @[RegSlices.scala 63:38 RegSlices.scala 66:41]
  assign fifo_h2c_cmd_io__in_bits_error = fifo_h2c_cmd_io_in_queue_io_downStream_bits_error; // @[RegSlices.scala 63:38 RegSlices.scala 66:41]
  assign fifo_h2c_cmd_io__in_bits_func = fifo_h2c_cmd_io_in_queue_io_downStream_bits_func; // @[RegSlices.scala 63:38 RegSlices.scala 66:41]
  assign fifo_h2c_cmd_io__in_bits_cidx = fifo_h2c_cmd_io_in_queue_io_downStream_bits_cidx; // @[RegSlices.scala 63:38 RegSlices.scala 66:41]
  assign fifo_h2c_cmd_io__in_bits_port_id = fifo_h2c_cmd_io_in_queue_io_downStream_bits_port_id; // @[RegSlices.scala 63:38 RegSlices.scala 66:41]
  assign fifo_h2c_cmd_io__in_bits_no_dma = fifo_h2c_cmd_io_in_queue_io_downStream_bits_no_dma; // @[RegSlices.scala 63:38 RegSlices.scala 66:41]
  assign fifo_h2c_cmd_io__out_ready = fifo_h2c_cmd_out_queue_io_upStream_ready; // @[RegSlices.scala 65:41]
  assign fifo_h2c_cmd_out_queue_clock = io_qdma_port_axi_aclk; // @[QDMADynamic.scala 47:53]
  assign fifo_h2c_cmd_out_queue_reset = ~io_qdma_port_axi_aresetn; // @[QDMADynamic.scala 58:64]
  assign fifo_h2c_cmd_out_queue_io_upStream_valid = fifo_h2c_cmd_io__out_valid; // @[RegSlices.scala 65:41]
  assign fifo_h2c_cmd_out_queue_io_upStream_bits_addr = fifo_h2c_cmd_io__out_bits_addr; // @[RegSlices.scala 65:41]
  assign fifo_h2c_cmd_out_queue_io_upStream_bits_len = fifo_h2c_cmd_io__out_bits_len; // @[RegSlices.scala 65:41]
  assign fifo_h2c_cmd_out_queue_io_upStream_bits_eop = fifo_h2c_cmd_io__out_bits_eop; // @[RegSlices.scala 65:41]
  assign fifo_h2c_cmd_out_queue_io_upStream_bits_sop = fifo_h2c_cmd_io__out_bits_sop; // @[RegSlices.scala 65:41]
  assign fifo_h2c_cmd_out_queue_io_upStream_bits_mrkr_req = fifo_h2c_cmd_io__out_bits_mrkr_req; // @[RegSlices.scala 65:41]
  assign fifo_h2c_cmd_out_queue_io_upStream_bits_sdi = fifo_h2c_cmd_io__out_bits_sdi; // @[RegSlices.scala 65:41]
  assign fifo_h2c_cmd_out_queue_io_upStream_bits_qid = fifo_h2c_cmd_io__out_bits_qid; // @[RegSlices.scala 65:41]
  assign fifo_h2c_cmd_out_queue_io_upStream_bits_error = fifo_h2c_cmd_io__out_bits_error; // @[RegSlices.scala 65:41]
  assign fifo_h2c_cmd_out_queue_io_upStream_bits_func = fifo_h2c_cmd_io__out_bits_func; // @[RegSlices.scala 65:41]
  assign fifo_h2c_cmd_out_queue_io_upStream_bits_cidx = fifo_h2c_cmd_io__out_bits_cidx; // @[RegSlices.scala 65:41]
  assign fifo_h2c_cmd_out_queue_io_upStream_bits_port_id = fifo_h2c_cmd_io__out_bits_port_id; // @[RegSlices.scala 65:41]
  assign fifo_h2c_cmd_out_queue_io_upStream_bits_no_dma = fifo_h2c_cmd_io__out_bits_no_dma; // @[RegSlices.scala 65:41]
  assign fifo_h2c_cmd_out_queue_io_downStream_ready = io_qdma_port_h2c_byp_in_st_rdy; // @[RegSlices.scala 63:38 QDMADynamic.scala 165:49]
  assign fifo_c2h_cmd_io_in_clk = io_user_clk; // @[XConverter.scala 62:33]
  assign fifo_c2h_cmd_io_out_clk = io_qdma_port_axi_aclk; // @[QDMADynamic.scala 47:53]
  assign fifo_c2h_cmd_io_rstn = io_user_arstn; // @[XConverter.scala 64:41]
  assign fifo_c2h_cmd_io_in_valid = boundary_split_io_cmd_out_valid; // @[QDMADynamic.scala 119:41]
  assign fifo_c2h_cmd_io_in_bits_addr = boundary_split_io_cmd_out_bits_addr; // @[QDMADynamic.scala 119:41]
  assign fifo_c2h_cmd_io_in_bits_qid = boundary_split_io_cmd_out_bits_qid; // @[QDMADynamic.scala 119:41]
  assign fifo_c2h_cmd_io_in_bits_error = boundary_split_io_cmd_out_bits_error; // @[QDMADynamic.scala 119:41]
  assign fifo_c2h_cmd_io_in_bits_func = boundary_split_io_cmd_out_bits_func; // @[QDMADynamic.scala 119:41]
  assign fifo_c2h_cmd_io_in_bits_port_id = boundary_split_io_cmd_out_bits_port_id; // @[QDMADynamic.scala 119:41]
  assign fifo_c2h_cmd_io_in_bits_pfch_tag = boundary_split_io_cmd_out_bits_pfch_tag; // @[QDMADynamic.scala 119:41]
  assign fifo_c2h_cmd_io_in_bits_len = boundary_split_io_cmd_out_bits_len; // @[QDMADynamic.scala 119:41]
  assign fifo_c2h_cmd_io_out_ready = fifo_c2h_cmd_out_queue_io_upStream_ready; // @[RegSlices.scala 65:41]
  assign fifo_c2h_cmd_out_queue_clock = io_qdma_port_axi_aclk; // @[QDMADynamic.scala 47:53]
  assign fifo_c2h_cmd_out_queue_reset = ~io_qdma_port_axi_aresetn; // @[QDMADynamic.scala 60:64]
  assign fifo_c2h_cmd_out_queue_io_upStream_valid = fifo_c2h_cmd_io_out_valid; // @[RegSlices.scala 65:41]
  assign fifo_c2h_cmd_out_queue_io_upStream_bits_addr = fifo_c2h_cmd_io_out_bits_addr; // @[RegSlices.scala 65:41]
  assign fifo_c2h_cmd_out_queue_io_upStream_bits_qid = fifo_c2h_cmd_io_out_bits_qid; // @[RegSlices.scala 65:41]
  assign fifo_c2h_cmd_out_queue_io_upStream_bits_error = fifo_c2h_cmd_io_out_bits_error; // @[RegSlices.scala 65:41]
  assign fifo_c2h_cmd_out_queue_io_upStream_bits_func = fifo_c2h_cmd_io_out_bits_func; // @[RegSlices.scala 65:41]
  assign fifo_c2h_cmd_out_queue_io_upStream_bits_port_id = fifo_c2h_cmd_io_out_bits_port_id; // @[RegSlices.scala 65:41]
  assign fifo_c2h_cmd_out_queue_io_upStream_bits_pfch_tag = fifo_c2h_cmd_io_out_bits_pfch_tag; // @[RegSlices.scala 65:41]
  assign fifo_c2h_cmd_out_queue_io_upStream_bits_len = fifo_c2h_cmd_io_out_bits_len; // @[RegSlices.scala 65:41]
  assign fifo_c2h_cmd_out_queue_io_downStream_ready = io_qdma_port_c2h_byp_in_st_csh_rdy; // @[RegSlices.scala 63:38 QDMADynamic.scala 175:57]
  assign check_c2h_clock = io_user_clk;
  assign check_c2h_reset = ~io_user_arstn; // @[QDMADynamic.scala 62:73]
  assign check_c2h_io_in_valid = check_c2h_io_in_queue_io_downStream_valid; // @[RegSlices.scala 63:38 RegSlices.scala 66:41]
  assign check_c2h_io_in_bits_addr = check_c2h_io_in_queue_io_downStream_bits_addr; // @[RegSlices.scala 63:38 RegSlices.scala 66:41]
  assign check_c2h_io_in_bits_qid = check_c2h_io_in_queue_io_downStream_bits_qid; // @[RegSlices.scala 63:38 RegSlices.scala 66:41]
  assign check_c2h_io_in_bits_error = check_c2h_io_in_queue_io_downStream_bits_error; // @[RegSlices.scala 63:38 RegSlices.scala 66:41]
  assign check_c2h_io_in_bits_func = check_c2h_io_in_queue_io_downStream_bits_func; // @[RegSlices.scala 63:38 RegSlices.scala 66:41]
  assign check_c2h_io_in_bits_port_id = check_c2h_io_in_queue_io_downStream_bits_port_id; // @[RegSlices.scala 63:38 RegSlices.scala 66:41]
  assign check_c2h_io_in_bits_pfch_tag = check_c2h_io_in_queue_io_downStream_bits_pfch_tag; // @[RegSlices.scala 63:38 RegSlices.scala 66:41]
  assign check_c2h_io_in_bits_len = check_c2h_io_in_queue_io_downStream_bits_len; // @[RegSlices.scala 63:38 RegSlices.scala 66:41]
  assign check_c2h_io_out_ready = tlb_io_c2h_in_queue_io_upStream_ready; // @[RegSlices.scala 65:41]
  assign check_c2h_io_in_queue_clock = io_user_clk;
  assign check_c2h_io_in_queue_reset = ~io_user_arstn; // @[QDMADynamic.scala 63:76]
  assign check_c2h_io_in_queue_io_upStream_valid = 1'h0; // @[RegSlices.scala 65:41]
  assign check_c2h_io_in_queue_io_upStream_bits_addr = 64'h0; // @[RegSlices.scala 65:41]
  assign check_c2h_io_in_queue_io_upStream_bits_qid = 11'h0; // @[RegSlices.scala 65:41]
  assign check_c2h_io_in_queue_io_upStream_bits_error = 1'h0; // @[RegSlices.scala 65:41]
  assign check_c2h_io_in_queue_io_upStream_bits_func = 8'h0; // @[RegSlices.scala 65:41]
  assign check_c2h_io_in_queue_io_upStream_bits_port_id = 3'h0; // @[RegSlices.scala 65:41]
  assign check_c2h_io_in_queue_io_upStream_bits_pfch_tag = 7'h0; // @[RegSlices.scala 65:41]
  assign check_c2h_io_in_queue_io_upStream_bits_len = 32'h0; // @[RegSlices.scala 65:41]
  assign check_c2h_io_in_queue_io_downStream_ready = check_c2h_io_in_ready; // @[RegSlices.scala 63:38 QDMADynamic.scala 63:41]
  assign check_h2c_clock = io_user_clk;
  assign check_h2c_reset = ~io_user_arstn; // @[QDMADynamic.scala 64:73]
  assign check_h2c_io_in_valid = check_h2c_io_in_queue_io_downStream_valid; // @[RegSlices.scala 63:38 RegSlices.scala 66:41]
  assign check_h2c_io_in_bits_addr = check_h2c_io_in_queue_io_downStream_bits_addr; // @[RegSlices.scala 63:38 RegSlices.scala 66:41]
  assign check_h2c_io_in_bits_len = check_h2c_io_in_queue_io_downStream_bits_len; // @[RegSlices.scala 63:38 RegSlices.scala 66:41]
  assign check_h2c_io_in_bits_eop = check_h2c_io_in_queue_io_downStream_bits_eop; // @[RegSlices.scala 63:38 RegSlices.scala 66:41]
  assign check_h2c_io_in_bits_sop = check_h2c_io_in_queue_io_downStream_bits_sop; // @[RegSlices.scala 63:38 RegSlices.scala 66:41]
  assign check_h2c_io_in_bits_mrkr_req = check_h2c_io_in_queue_io_downStream_bits_mrkr_req; // @[RegSlices.scala 63:38 RegSlices.scala 66:41]
  assign check_h2c_io_in_bits_sdi = check_h2c_io_in_queue_io_downStream_bits_sdi; // @[RegSlices.scala 63:38 RegSlices.scala 66:41]
  assign check_h2c_io_in_bits_qid = check_h2c_io_in_queue_io_downStream_bits_qid; // @[RegSlices.scala 63:38 RegSlices.scala 66:41]
  assign check_h2c_io_in_bits_error = check_h2c_io_in_queue_io_downStream_bits_error; // @[RegSlices.scala 63:38 RegSlices.scala 66:41]
  assign check_h2c_io_in_bits_func = check_h2c_io_in_queue_io_downStream_bits_func; // @[RegSlices.scala 63:38 RegSlices.scala 66:41]
  assign check_h2c_io_in_bits_cidx = check_h2c_io_in_queue_io_downStream_bits_cidx; // @[RegSlices.scala 63:38 RegSlices.scala 66:41]
  assign check_h2c_io_in_bits_port_id = check_h2c_io_in_queue_io_downStream_bits_port_id; // @[RegSlices.scala 63:38 RegSlices.scala 66:41]
  assign check_h2c_io_in_bits_no_dma = check_h2c_io_in_queue_io_downStream_bits_no_dma; // @[RegSlices.scala 63:38 RegSlices.scala 66:41]
  assign check_h2c_io_out_ready = tlb_io_h2c_in_queue_io_upStream_ready; // @[RegSlices.scala 65:41]
  assign check_h2c_io_in_queue_clock = io_user_clk;
  assign check_h2c_io_in_queue_reset = ~io_user_arstn; // @[QDMADynamic.scala 65:76]
  assign check_h2c_io_in_queue_io_upStream_valid = io_h2c_cmd_valid; // @[RegSlices.scala 65:41]
  assign check_h2c_io_in_queue_io_upStream_bits_addr = io_h2c_cmd_bits_addr; // @[RegSlices.scala 65:41]
  assign check_h2c_io_in_queue_io_upStream_bits_len = io_h2c_cmd_bits_len; // @[RegSlices.scala 65:41]
  assign check_h2c_io_in_queue_io_upStream_bits_eop = 1'h1; // @[RegSlices.scala 65:41]
  assign check_h2c_io_in_queue_io_upStream_bits_sop = 1'h1; // @[RegSlices.scala 65:41]
  assign check_h2c_io_in_queue_io_upStream_bits_mrkr_req = 1'h0; // @[RegSlices.scala 65:41]
  assign check_h2c_io_in_queue_io_upStream_bits_sdi = 1'h0; // @[RegSlices.scala 65:41]
  assign check_h2c_io_in_queue_io_upStream_bits_qid = 11'h0; // @[RegSlices.scala 65:41]
  assign check_h2c_io_in_queue_io_upStream_bits_error = 1'h0; // @[RegSlices.scala 65:41]
  assign check_h2c_io_in_queue_io_upStream_bits_func = 8'h0; // @[RegSlices.scala 65:41]
  assign check_h2c_io_in_queue_io_upStream_bits_cidx = 16'h0; // @[RegSlices.scala 65:41]
  assign check_h2c_io_in_queue_io_upStream_bits_port_id = 3'h0; // @[RegSlices.scala 65:41]
  assign check_h2c_io_in_queue_io_upStream_bits_no_dma = 1'h0; // @[RegSlices.scala 65:41]
  assign check_h2c_io_in_queue_io_downStream_ready = check_h2c_io_in_ready; // @[RegSlices.scala 63:38 QDMADynamic.scala 65:41]
  assign tlb_clock = io_user_clk;
  assign tlb_reset = ~io_user_arstn; // @[QDMADynamic.scala 67:49]
  assign tlb_io__wr_tlb_valid = wr_tlb_valid_REG_1; // @[QDMADynamic.scala 74:39 QDMADynamic.scala 81:33]
  assign tlb_io__wr_tlb_bits_vaddr_high = io_reg_control_9; // @[QDMADynamic.scala 74:39 QDMADynamic.scala 78:33]
  assign tlb_io__wr_tlb_bits_vaddr_low = io_reg_control_8; // @[QDMADynamic.scala 74:39 QDMADynamic.scala 79:33]
  assign tlb_io__wr_tlb_bits_paddr_high = io_reg_control_11; // @[QDMADynamic.scala 74:39 QDMADynamic.scala 76:33]
  assign tlb_io__wr_tlb_bits_paddr_low = io_reg_control_10; // @[QDMADynamic.scala 74:39 QDMADynamic.scala 77:33]
  assign tlb_io__wr_tlb_bits_is_base = io_reg_control_12[0]; // @[QDMADynamic.scala 75:62]
  assign tlb_io__h2c_in_valid = tlb_io_h2c_in_queue_io_downStream_valid; // @[RegSlices.scala 63:38 RegSlices.scala 66:41]
  assign tlb_io__h2c_in_bits_addr = tlb_io_h2c_in_queue_io_downStream_bits_addr; // @[RegSlices.scala 63:38 RegSlices.scala 66:41]
  assign tlb_io__h2c_in_bits_len = tlb_io_h2c_in_queue_io_downStream_bits_len; // @[RegSlices.scala 63:38 RegSlices.scala 66:41]
  assign tlb_io__h2c_in_bits_eop = tlb_io_h2c_in_queue_io_downStream_bits_eop; // @[RegSlices.scala 63:38 RegSlices.scala 66:41]
  assign tlb_io__h2c_in_bits_sop = tlb_io_h2c_in_queue_io_downStream_bits_sop; // @[RegSlices.scala 63:38 RegSlices.scala 66:41]
  assign tlb_io__h2c_in_bits_mrkr_req = tlb_io_h2c_in_queue_io_downStream_bits_mrkr_req; // @[RegSlices.scala 63:38 RegSlices.scala 66:41]
  assign tlb_io__h2c_in_bits_sdi = tlb_io_h2c_in_queue_io_downStream_bits_sdi; // @[RegSlices.scala 63:38 RegSlices.scala 66:41]
  assign tlb_io__h2c_in_bits_qid = tlb_io_h2c_in_queue_io_downStream_bits_qid; // @[RegSlices.scala 63:38 RegSlices.scala 66:41]
  assign tlb_io__h2c_in_bits_error = tlb_io_h2c_in_queue_io_downStream_bits_error; // @[RegSlices.scala 63:38 RegSlices.scala 66:41]
  assign tlb_io__h2c_in_bits_func = tlb_io_h2c_in_queue_io_downStream_bits_func; // @[RegSlices.scala 63:38 RegSlices.scala 66:41]
  assign tlb_io__h2c_in_bits_cidx = tlb_io_h2c_in_queue_io_downStream_bits_cidx; // @[RegSlices.scala 63:38 RegSlices.scala 66:41]
  assign tlb_io__h2c_in_bits_port_id = tlb_io_h2c_in_queue_io_downStream_bits_port_id; // @[RegSlices.scala 63:38 RegSlices.scala 66:41]
  assign tlb_io__h2c_in_bits_no_dma = tlb_io_h2c_in_queue_io_downStream_bits_no_dma; // @[RegSlices.scala 63:38 RegSlices.scala 66:41]
  assign tlb_io__c2h_in_valid = tlb_io_c2h_in_queue_io_downStream_valid; // @[RegSlices.scala 63:38 RegSlices.scala 66:41]
  assign tlb_io__c2h_in_bits_addr = tlb_io_c2h_in_queue_io_downStream_bits_addr; // @[RegSlices.scala 63:38 RegSlices.scala 66:41]
  assign tlb_io__c2h_in_bits_qid = tlb_io_c2h_in_queue_io_downStream_bits_qid; // @[RegSlices.scala 63:38 RegSlices.scala 66:41]
  assign tlb_io__c2h_in_bits_error = tlb_io_c2h_in_queue_io_downStream_bits_error; // @[RegSlices.scala 63:38 RegSlices.scala 66:41]
  assign tlb_io__c2h_in_bits_func = tlb_io_c2h_in_queue_io_downStream_bits_func; // @[RegSlices.scala 63:38 RegSlices.scala 66:41]
  assign tlb_io__c2h_in_bits_port_id = tlb_io_c2h_in_queue_io_downStream_bits_port_id; // @[RegSlices.scala 63:38 RegSlices.scala 66:41]
  assign tlb_io__c2h_in_bits_pfch_tag = tlb_io_c2h_in_queue_io_downStream_bits_pfch_tag; // @[RegSlices.scala 63:38 RegSlices.scala 66:41]
  assign tlb_io__c2h_in_bits_len = tlb_io_c2h_in_queue_io_downStream_bits_len; // @[RegSlices.scala 63:38 RegSlices.scala 66:41]
  assign tlb_io__h2c_out_ready = fifo_h2c_cmd_io_in_queue_io_upStream_ready; // @[RegSlices.scala 65:41]
  assign tlb_io__c2h_out_ready = boundary_split_io_cmd_in_ready; // @[QDMADynamic.scala 117:34]
  assign tlb_io_h2c_in_queue_clock = io_user_clk;
  assign tlb_io_h2c_in_queue_reset = ~io_user_arstn; // @[QDMADynamic.scala 69:68]
  assign tlb_io_h2c_in_queue_io_upStream_valid = check_h2c_io_out_valid; // @[RegSlices.scala 65:41]
  assign tlb_io_h2c_in_queue_io_upStream_bits_addr = check_h2c_io_out_bits_addr; // @[RegSlices.scala 65:41]
  assign tlb_io_h2c_in_queue_io_upStream_bits_len = check_h2c_io_out_bits_len; // @[RegSlices.scala 65:41]
  assign tlb_io_h2c_in_queue_io_upStream_bits_eop = check_h2c_io_out_bits_eop; // @[RegSlices.scala 65:41]
  assign tlb_io_h2c_in_queue_io_upStream_bits_sop = check_h2c_io_out_bits_sop; // @[RegSlices.scala 65:41]
  assign tlb_io_h2c_in_queue_io_upStream_bits_mrkr_req = check_h2c_io_out_bits_mrkr_req; // @[RegSlices.scala 65:41]
  assign tlb_io_h2c_in_queue_io_upStream_bits_sdi = check_h2c_io_out_bits_sdi; // @[RegSlices.scala 65:41]
  assign tlb_io_h2c_in_queue_io_upStream_bits_qid = check_h2c_io_out_bits_qid; // @[RegSlices.scala 65:41]
  assign tlb_io_h2c_in_queue_io_upStream_bits_error = check_h2c_io_out_bits_error; // @[RegSlices.scala 65:41]
  assign tlb_io_h2c_in_queue_io_upStream_bits_func = check_h2c_io_out_bits_func; // @[RegSlices.scala 65:41]
  assign tlb_io_h2c_in_queue_io_upStream_bits_cidx = check_h2c_io_out_bits_cidx; // @[RegSlices.scala 65:41]
  assign tlb_io_h2c_in_queue_io_upStream_bits_port_id = check_h2c_io_out_bits_port_id; // @[RegSlices.scala 65:41]
  assign tlb_io_h2c_in_queue_io_upStream_bits_no_dma = check_h2c_io_out_bits_no_dma; // @[RegSlices.scala 65:41]
  assign tlb_io_h2c_in_queue_io_downStream_ready = tlb_io__h2c_in_ready; // @[RegSlices.scala 63:38 QDMADynamic.scala 69:33]
  assign tlb_io_c2h_in_queue_clock = io_user_clk;
  assign tlb_io_c2h_in_queue_reset = ~io_user_arstn; // @[QDMADynamic.scala 70:68]
  assign tlb_io_c2h_in_queue_io_upStream_valid = check_c2h_io_out_valid; // @[RegSlices.scala 65:41]
  assign tlb_io_c2h_in_queue_io_upStream_bits_addr = check_c2h_io_out_bits_addr; // @[RegSlices.scala 65:41]
  assign tlb_io_c2h_in_queue_io_upStream_bits_qid = check_c2h_io_out_bits_qid; // @[RegSlices.scala 65:41]
  assign tlb_io_c2h_in_queue_io_upStream_bits_error = check_c2h_io_out_bits_error; // @[RegSlices.scala 65:41]
  assign tlb_io_c2h_in_queue_io_upStream_bits_func = check_c2h_io_out_bits_func; // @[RegSlices.scala 65:41]
  assign tlb_io_c2h_in_queue_io_upStream_bits_port_id = check_c2h_io_out_bits_port_id; // @[RegSlices.scala 65:41]
  assign tlb_io_c2h_in_queue_io_upStream_bits_pfch_tag = check_c2h_io_out_bits_pfch_tag; // @[RegSlices.scala 65:41]
  assign tlb_io_c2h_in_queue_io_upStream_bits_len = check_c2h_io_out_bits_len; // @[RegSlices.scala 65:41]
  assign tlb_io_c2h_in_queue_io_downStream_ready = tlb_io__c2h_in_ready; // @[RegSlices.scala 63:38 QDMADynamic.scala 70:33]
  assign fifo_h2c_cmd_io_in_queue_clock = io_user_clk;
  assign fifo_h2c_cmd_io_in_queue_reset = ~io_user_arstn; // @[QDMADynamic.scala 71:68]
  assign fifo_h2c_cmd_io_in_queue_io_upStream_valid = tlb_io__h2c_out_valid; // @[RegSlices.scala 65:41]
  assign fifo_h2c_cmd_io_in_queue_io_upStream_bits_addr = tlb_io__h2c_out_bits_addr; // @[RegSlices.scala 65:41]
  assign fifo_h2c_cmd_io_in_queue_io_upStream_bits_len = tlb_io__h2c_out_bits_len; // @[RegSlices.scala 65:41]
  assign fifo_h2c_cmd_io_in_queue_io_upStream_bits_eop = tlb_io__h2c_out_bits_eop; // @[RegSlices.scala 65:41]
  assign fifo_h2c_cmd_io_in_queue_io_upStream_bits_sop = tlb_io__h2c_out_bits_sop; // @[RegSlices.scala 65:41]
  assign fifo_h2c_cmd_io_in_queue_io_upStream_bits_mrkr_req = tlb_io__h2c_out_bits_mrkr_req; // @[RegSlices.scala 65:41]
  assign fifo_h2c_cmd_io_in_queue_io_upStream_bits_sdi = tlb_io__h2c_out_bits_sdi; // @[RegSlices.scala 65:41]
  assign fifo_h2c_cmd_io_in_queue_io_upStream_bits_qid = tlb_io__h2c_out_bits_qid; // @[RegSlices.scala 65:41]
  assign fifo_h2c_cmd_io_in_queue_io_upStream_bits_error = tlb_io__h2c_out_bits_error; // @[RegSlices.scala 65:41]
  assign fifo_h2c_cmd_io_in_queue_io_upStream_bits_func = tlb_io__h2c_out_bits_func; // @[RegSlices.scala 65:41]
  assign fifo_h2c_cmd_io_in_queue_io_upStream_bits_cidx = tlb_io__h2c_out_bits_cidx; // @[RegSlices.scala 65:41]
  assign fifo_h2c_cmd_io_in_queue_io_upStream_bits_port_id = tlb_io__h2c_out_bits_port_id; // @[RegSlices.scala 65:41]
  assign fifo_h2c_cmd_io_in_queue_io_upStream_bits_no_dma = tlb_io__h2c_out_bits_no_dma; // @[RegSlices.scala 65:41]
  assign fifo_h2c_cmd_io_in_queue_io_downStream_ready = fifo_h2c_cmd_io__in_ready; // @[RegSlices.scala 63:38 QDMADynamic.scala 71:33]
  assign axil2reg_clock = io_user_clk;
  assign axil2reg_reset = ~io_user_arstn; // @[QDMADynamic.scala 86:54]
  assign axil2reg_io_axi_aw_valid = axil2reg_io_axi_cvt_aw_io_out_valid; // @[XConverter.scala 22:39 XConverter.scala 41:33]
  assign axil2reg_io_axi_aw_bits_addr = axil2reg_io_axi_cvt_aw_io_out_bits_addr; // @[XConverter.scala 22:39 XConverter.scala 41:33]
  assign axil2reg_io_axi_ar_valid = axil2reg_io_axi_cvt_ar_io_out_valid; // @[XConverter.scala 22:39 XConverter.scala 42:33]
  assign axil2reg_io_axi_ar_bits_addr = axil2reg_io_axi_cvt_ar_io_out_bits_addr; // @[XConverter.scala 22:39 XConverter.scala 42:33]
  assign axil2reg_io_axi_w_valid = axil2reg_io_axi_cvt_w_io_out_valid; // @[XConverter.scala 22:39 XConverter.scala 43:33]
  assign axil2reg_io_axi_w_bits_data = axil2reg_io_axi_cvt_w_io_out_bits_data; // @[XConverter.scala 22:39 XConverter.scala 43:33]
  assign axil2reg_io_axi_r_ready = axil2reg_io_axi_cvt_r_io_in_ready; // @[XConverter.scala 22:39 XConverter.scala 44:41]
  assign axil2reg_io_reg_status_300 = io_reg_status_300; // @[QDMADynamic.scala 88:33]
  assign axil2reg_io_reg_status_400 = io_reg_status_400; // @[QDMADynamic.scala 88:33]
  assign axil2reg_io_reg_status_401 = io_reg_status_401; // @[QDMADynamic.scala 88:33]
  assign axil2reg_io_reg_status_402 = io_reg_status_402; // @[QDMADynamic.scala 88:33]
  assign axil2reg_io_reg_status_403 = io_reg_status_403; // @[QDMADynamic.scala 88:33]
  assign axil2reg_io_reg_status_404 = io_reg_status_404; // @[QDMADynamic.scala 88:33]
  assign axil2reg_io_reg_status_405 = io_reg_status_405; // @[QDMADynamic.scala 88:33]
  assign axil2reg_io_reg_status_406 = io_reg_status_406; // @[QDMADynamic.scala 88:33]
  assign axil2reg_io_reg_status_407 = io_reg_status_407; // @[QDMADynamic.scala 88:33]
  assign axil2reg_io_reg_status_408 = io_reg_status_408; // @[QDMADynamic.scala 88:33]
  assign axil2reg_io_reg_status_409 = io_reg_status_409; // @[QDMADynamic.scala 88:33]
  assign axil2reg_io_reg_status_410 = io_reg_status_410; // @[QDMADynamic.scala 88:33]
  assign axil2reg_io_reg_status_411 = io_reg_status_411; // @[QDMADynamic.scala 88:33]
  assign axil2reg_io_reg_status_412 = io_reg_status_412; // @[QDMADynamic.scala 88:33]
  assign axil2reg_io_reg_status_413 = io_reg_status_413; // @[QDMADynamic.scala 88:33]
  assign axil2reg_io_reg_status_414 = io_reg_status_414; // @[QDMADynamic.scala 88:33]
  assign io_axib_cvt_aw_io_in_clk = io_qdma_port_axi_aclk; // @[QDMADynamic.scala 47:53]
  assign io_axib_cvt_aw_io_out_clk = io_user_clk; // @[XConverter.scala 63:33]
  assign io_axib_cvt_aw_io_rstn = io_qdma_port_axi_aresetn; // @[QDMADynamic.scala 48:51]
  assign io_axib_cvt_aw_io_in_valid = io_qdma_port_m_axib_awvalid; // @[QDMADynamic.scala 92:24 QDMADynamic.scala 212:65]
  assign io_axib_cvt_aw_io_in_bits_addr = io_qdma_port_m_axib_awaddr; // @[QDMADynamic.scala 92:24 QDMADynamic.scala 205:65]
  assign io_axib_cvt_aw_io_in_bits_burst = io_qdma_port_m_axib_awburst; // @[QDMADynamic.scala 92:24 QDMADynamic.scala 208:65]
  assign io_axib_cvt_aw_io_in_bits_cache = io_qdma_port_m_axib_awcache; // @[QDMADynamic.scala 92:24 QDMADynamic.scala 211:65]
  assign io_axib_cvt_aw_io_in_bits_id = io_qdma_port_m_axib_awid; // @[QDMADynamic.scala 92:24 QDMADynamic.scala 204:65]
  assign io_axib_cvt_aw_io_in_bits_len = io_qdma_port_m_axib_awlen; // @[QDMADynamic.scala 92:24 QDMADynamic.scala 206:65]
  assign io_axib_cvt_aw_io_in_bits_lock = io_qdma_port_m_axib_awlock; // @[QDMADynamic.scala 92:24 QDMADynamic.scala 210:65]
  assign io_axib_cvt_aw_io_in_bits_prot = io_qdma_port_m_axib_awprot; // @[QDMADynamic.scala 92:24 QDMADynamic.scala 209:65]
  assign io_axib_cvt_aw_io_in_bits_size = io_qdma_port_m_axib_awsize; // @[QDMADynamic.scala 92:24 QDMADynamic.scala 207:65]
  assign io_axib_cvt_aw_io_out_ready = io_axib_aw_ready; // @[XConverter.scala 22:39 QDMADynamic.scala 96:17]
  assign io_axib_cvt_ar_io_in_clk = io_qdma_port_axi_aclk; // @[QDMADynamic.scala 47:53]
  assign io_axib_cvt_ar_io_out_clk = io_user_clk; // @[XConverter.scala 63:33]
  assign io_axib_cvt_ar_io_rstn = io_qdma_port_axi_aresetn; // @[QDMADynamic.scala 48:51]
  assign io_axib_cvt_ar_io_in_valid = io_qdma_port_m_axib_arvalid; // @[QDMADynamic.scala 92:24 QDMADynamic.scala 234:65]
  assign io_axib_cvt_ar_io_in_bits_addr = io_qdma_port_m_axib_araddr; // @[QDMADynamic.scala 92:24 QDMADynamic.scala 227:65]
  assign io_axib_cvt_ar_io_in_bits_burst = io_qdma_port_m_axib_arburst; // @[QDMADynamic.scala 92:24 QDMADynamic.scala 230:65]
  assign io_axib_cvt_ar_io_in_bits_cache = io_qdma_port_m_axib_arcache; // @[QDMADynamic.scala 92:24 QDMADynamic.scala 233:65]
  assign io_axib_cvt_ar_io_in_bits_id = io_qdma_port_m_axib_arid; // @[QDMADynamic.scala 92:24 QDMADynamic.scala 226:65]
  assign io_axib_cvt_ar_io_in_bits_len = io_qdma_port_m_axib_arlen; // @[QDMADynamic.scala 92:24 QDMADynamic.scala 228:65]
  assign io_axib_cvt_ar_io_in_bits_lock = io_qdma_port_m_axib_arlock; // @[QDMADynamic.scala 92:24 QDMADynamic.scala 232:65]
  assign io_axib_cvt_ar_io_in_bits_prot = io_qdma_port_m_axib_arprot; // @[QDMADynamic.scala 92:24 QDMADynamic.scala 231:65]
  assign io_axib_cvt_ar_io_in_bits_size = io_qdma_port_m_axib_arsize; // @[QDMADynamic.scala 92:24 QDMADynamic.scala 229:65]
  assign io_axib_cvt_ar_io_out_ready = 1'h1; // @[XConverter.scala 22:39 QDMADynamic.scala 96:17]
  assign io_axib_cvt_w_io_in_clk = io_qdma_port_axi_aclk; // @[QDMADynamic.scala 47:53]
  assign io_axib_cvt_w_io_out_clk = io_user_clk; // @[XConverter.scala 63:33]
  assign io_axib_cvt_w_io_rstn = io_qdma_port_axi_aresetn; // @[QDMADynamic.scala 48:51]
  assign io_axib_cvt_w_io_in_valid = io_qdma_port_m_axib_wvalid; // @[QDMADynamic.scala 92:24 QDMADynamic.scala 218:65]
  assign io_axib_cvt_w_io_in_bits_data = io_qdma_port_m_axib_wdata; // @[QDMADynamic.scala 92:24 QDMADynamic.scala 215:65]
  assign io_axib_cvt_w_io_in_bits_last = io_qdma_port_m_axib_wlast; // @[QDMADynamic.scala 92:24 QDMADynamic.scala 217:65]
  assign io_axib_cvt_w_io_in_bits_strb = io_qdma_port_m_axib_wstrb; // @[QDMADynamic.scala 92:24 QDMADynamic.scala 216:65]
  assign io_axib_cvt_w_io_out_ready = io_axib_w_ready; // @[XConverter.scala 22:39 QDMADynamic.scala 96:17]
  assign io_axib_cvt_r_io_in_clk = io_user_clk; // @[XConverter.scala 62:33]
  assign io_axib_cvt_r_io_out_clk = io_qdma_port_axi_aclk; // @[QDMADynamic.scala 47:53]
  assign io_axib_cvt_r_io_rstn = io_user_arstn; // @[XConverter.scala 64:41]
  assign io_axib_cvt_r_io_in_bits_data = io_axib_r_bits_data; // @[XConverter.scala 22:39 QDMADynamic.scala 96:17]
  assign io_axib_cvt_r_io_out_ready = io_qdma_port_m_axib_rready; // @[QDMADynamic.scala 92:24 QDMADynamic.scala 242:65]
  assign io_axib_cvt_b_io_in_clk = io_user_clk; // @[XConverter.scala 62:33]
  assign io_axib_cvt_b_io_out_clk = io_qdma_port_axi_aclk; // @[QDMADynamic.scala 47:53]
  assign io_axib_cvt_b_io_rstn = io_user_arstn; // @[XConverter.scala 64:41]
  assign io_axib_cvt_b_io_out_ready = io_qdma_port_m_axib_bready; // @[QDMADynamic.scala 92:24 QDMADynamic.scala 224:65]
  assign axil2reg_io_axi_cvt_aw_io_in_clk = io_qdma_port_axi_aclk; // @[QDMADynamic.scala 47:53]
  assign axil2reg_io_axi_cvt_aw_io_out_clk = io_user_clk; // @[XConverter.scala 63:33]
  assign axil2reg_io_axi_cvt_aw_io_rstn = io_qdma_port_axi_aresetn; // @[QDMADynamic.scala 48:51]
  assign axil2reg_io_axi_cvt_aw_io_in_valid = io_qdma_port_m_axil_awvalid; // @[QDMADynamic.scala 107:24 QDMADynamic.scala 245:65]
  assign axil2reg_io_axi_cvt_aw_io_in_bits_addr = io_qdma_port_m_axil_awaddr; // @[QDMADynamic.scala 107:24 QDMADynamic.scala 244:65]
  assign axil2reg_io_axi_cvt_aw_io_out_ready = axil2reg_io_axi_aw_ready; // @[XConverter.scala 22:39 QDMADynamic.scala 113:25]
  assign axil2reg_io_axi_cvt_ar_io_in_clk = io_qdma_port_axi_aclk; // @[QDMADynamic.scala 47:53]
  assign axil2reg_io_axi_cvt_ar_io_out_clk = io_user_clk; // @[XConverter.scala 63:33]
  assign axil2reg_io_axi_cvt_ar_io_rstn = io_qdma_port_axi_aresetn; // @[QDMADynamic.scala 48:51]
  assign axil2reg_io_axi_cvt_ar_io_in_valid = io_qdma_port_m_axil_arvalid; // @[QDMADynamic.scala 107:24 QDMADynamic.scala 258:65]
  assign axil2reg_io_axi_cvt_ar_io_in_bits_addr = io_qdma_port_m_axil_araddr; // @[QDMADynamic.scala 107:24 QDMADynamic.scala 257:65]
  assign axil2reg_io_axi_cvt_ar_io_out_ready = axil2reg_io_axi_ar_ready; // @[XConverter.scala 22:39 QDMADynamic.scala 113:25]
  assign axil2reg_io_axi_cvt_w_io_in_clk = io_qdma_port_axi_aclk; // @[QDMADynamic.scala 47:53]
  assign axil2reg_io_axi_cvt_w_io_out_clk = io_user_clk; // @[XConverter.scala 63:33]
  assign axil2reg_io_axi_cvt_w_io_rstn = io_qdma_port_axi_aresetn; // @[QDMADynamic.scala 48:51]
  assign axil2reg_io_axi_cvt_w_io_in_valid = io_qdma_port_m_axil_wvalid; // @[QDMADynamic.scala 107:24 QDMADynamic.scala 250:65]
  assign axil2reg_io_axi_cvt_w_io_in_bits_data = io_qdma_port_m_axil_wdata; // @[QDMADynamic.scala 107:24 QDMADynamic.scala 248:65]
  assign axil2reg_io_axi_cvt_w_io_in_bits_strb = io_qdma_port_m_axil_wstrb; // @[QDMADynamic.scala 107:24 QDMADynamic.scala 249:65]
  assign axil2reg_io_axi_cvt_w_io_out_ready = axil2reg_io_axi_w_ready; // @[XConverter.scala 22:39 QDMADynamic.scala 113:25]
  assign axil2reg_io_axi_cvt_r_io_in_clk = io_user_clk; // @[XConverter.scala 62:33]
  assign axil2reg_io_axi_cvt_r_io_out_clk = io_qdma_port_axi_aclk; // @[QDMADynamic.scala 47:53]
  assign axil2reg_io_axi_cvt_r_io_rstn = io_user_arstn; // @[XConverter.scala 64:41]
  assign axil2reg_io_axi_cvt_r_io_in_valid = axil2reg_io_axi_r_valid; // @[XConverter.scala 22:39 QDMADynamic.scala 113:25]
  assign axil2reg_io_axi_cvt_r_io_in_bits_data = axil2reg_io_axi_r_bits_data; // @[XConverter.scala 22:39 QDMADynamic.scala 113:25]
  assign axil2reg_io_axi_cvt_r_io_out_ready = io_qdma_port_m_axil_rready; // @[QDMADynamic.scala 107:24 QDMADynamic.scala 264:65]
  assign axil2reg_io_axi_cvt_b_io_in_clk = io_user_clk; // @[XConverter.scala 62:33]
  assign axil2reg_io_axi_cvt_b_io_out_clk = io_qdma_port_axi_aclk; // @[QDMADynamic.scala 47:53]
  assign axil2reg_io_axi_cvt_b_io_rstn = io_user_arstn; // @[XConverter.scala 64:41]
  assign axil2reg_io_axi_cvt_b_io_out_ready = io_qdma_port_m_axil_bready; // @[QDMADynamic.scala 107:24 QDMADynamic.scala 255:65]
  assign boundary_split_clock = io_user_clk;
  assign boundary_split_reset = ~io_user_arstn; // @[QDMADynamic.scala 116:60]
  assign boundary_split_io_cmd_in_valid = tlb_io__c2h_out_valid; // @[QDMADynamic.scala 117:34]
  assign boundary_split_io_cmd_in_bits_addr = tlb_io__c2h_out_bits_addr; // @[QDMADynamic.scala 117:34]
  assign boundary_split_io_cmd_in_bits_qid = tlb_io__c2h_out_bits_qid; // @[QDMADynamic.scala 117:34]
  assign boundary_split_io_cmd_in_bits_error = tlb_io__c2h_out_bits_error; // @[QDMADynamic.scala 117:34]
  assign boundary_split_io_cmd_in_bits_func = tlb_io__c2h_out_bits_func; // @[QDMADynamic.scala 117:34]
  assign boundary_split_io_cmd_in_bits_port_id = tlb_io__c2h_out_bits_port_id; // @[QDMADynamic.scala 117:34]
  assign boundary_split_io_cmd_in_bits_pfch_tag = tlb_io__c2h_out_bits_pfch_tag; // @[QDMADynamic.scala 117:34]
  assign boundary_split_io_cmd_in_bits_len = tlb_io__c2h_out_bits_len; // @[QDMADynamic.scala 117:34]
  assign boundary_split_io_data_out_ready = fifo_c2h_data_io__in_ready; // @[QDMADynamic.scala 120:41]
  assign boundary_split_io_cmd_out_ready = fifo_c2h_cmd_io_in_ready; // @[QDMADynamic.scala 119:41]
  always @(posedge io_user_clk) begin
    wr_tlb_valid_REG <= io_reg_control_13[0]; // @[QDMADynamic.scala 81:118]
    wr_tlb_valid_REG_1 <= ~wr_tlb_valid_REG & io_reg_control_13[0]; // @[QDMADynamic.scala 81:123]
    if (_T_6) begin // @[Collector.scala 169:42]
      counter <= 32'h0; // @[Collector.scala 169:42]
    end
    if (_T_6) begin // @[Collector.scala 169:42]
      counter_1 <= 32'h0; // @[Collector.scala 169:42]
    end else if (_T_8) begin // @[Collector.scala 170:34]
      counter_1 <= _counter_T_3; // @[Collector.scala 171:41]
    end
    if (_T_6) begin // @[Collector.scala 169:42]
      counter_2 <= 32'h0; // @[Collector.scala 169:42]
    end
    if (_T_6) begin // @[Collector.scala 169:42]
      counter_3 <= 32'h0; // @[Collector.scala 169:42]
    end else if (io_h2c_data_valid) begin // @[Collector.scala 170:34]
      counter_3 <= _counter_T_7; // @[Collector.scala 171:41]
    end
  end
  always @(posedge io_qdma_port_axi_aclk) begin
    if (_T_12) begin // @[Collector.scala 169:42]
      counter_4 <= 32'h0; // @[Collector.scala 169:42]
    end else if (_T_13) begin // @[Collector.scala 170:34]
      counter_4 <= _counter_T_9; // @[Collector.scala 171:41]
    end
    if (_T_12) begin // @[Collector.scala 169:42]
      counter_5 <= 32'h0; // @[Collector.scala 169:42]
    end else if (_T_14) begin // @[Collector.scala 170:34]
      counter_5 <= _counter_T_11; // @[Collector.scala 171:41]
    end
    if (_T_12) begin // @[Collector.scala 169:42]
      counter_6 <= 32'h0; // @[Collector.scala 169:42]
    end else if (_T_15) begin // @[Collector.scala 170:34]
      counter_6 <= _counter_T_13; // @[Collector.scala 171:41]
    end
    if (_T_12) begin // @[Collector.scala 169:42]
      counter_7 <= 32'h0; // @[Collector.scala 169:42]
    end else if (_T_16) begin // @[Collector.scala 170:34]
      counter_7 <= _counter_T_15; // @[Collector.scala 171:41]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  wr_tlb_valid_REG = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  wr_tlb_valid_REG_1 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  counter = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  counter_1 = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  counter_2 = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  counter_3 = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  counter_4 = _RAND_6[31:0];
  _RAND_7 = {1{`RANDOM}};
  counter_5 = _RAND_7[31:0];
  _RAND_8 = {1{`RANDOM}};
  counter_6 = _RAND_8[31:0];
  _RAND_9 = {1{`RANDOM}};
  counter_7 = _RAND_9[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Queue_4(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input  [9:0]  io_enq_bits_class_id,
  input  [63:0] io_enq_bits_host_base_addr,
  input         io_deq_ready,
  output        io_deq_valid,
  output [9:0]  io_deq_bits_class_id,
  output [63:0] io_deq_bits_host_base_addr
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
  reg [63:0] _RAND_1;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
`endif // RANDOMIZE_REG_INIT
  reg [9:0] ram_class_id [0:7]; // @[Decoupled.scala 218:16]
  wire [9:0] ram_class_id_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16]
  wire [2:0] ram_class_id_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16]
  wire [9:0] ram_class_id_MPORT_data; // @[Decoupled.scala 218:16]
  wire [2:0] ram_class_id_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_class_id_MPORT_mask; // @[Decoupled.scala 218:16]
  wire  ram_class_id_MPORT_en; // @[Decoupled.scala 218:16]
  reg [63:0] ram_host_base_addr [0:7]; // @[Decoupled.scala 218:16]
  wire [63:0] ram_host_base_addr_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16]
  wire [2:0] ram_host_base_addr_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16]
  wire [63:0] ram_host_base_addr_MPORT_data; // @[Decoupled.scala 218:16]
  wire [2:0] ram_host_base_addr_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_host_base_addr_MPORT_mask; // @[Decoupled.scala 218:16]
  wire  ram_host_base_addr_MPORT_en; // @[Decoupled.scala 218:16]
  reg [2:0] enq_ptr_value; // @[Counter.scala 60:40]
  reg [2:0] deq_ptr_value; // @[Counter.scala 60:40]
  reg  maybe_full; // @[Decoupled.scala 221:27]
  wire  ptr_match = enq_ptr_value == deq_ptr_value; // @[Decoupled.scala 223:33]
  wire  empty = ptr_match & ~maybe_full; // @[Decoupled.scala 224:25]
  wire  full = ptr_match & maybe_full; // @[Decoupled.scala 225:24]
  wire  do_enq = io_enq_ready & io_enq_valid; // @[Decoupled.scala 40:37]
  wire  do_deq = io_deq_ready & io_deq_valid; // @[Decoupled.scala 40:37]
  wire [2:0] _value_T_1 = enq_ptr_value + 3'h1; // @[Counter.scala 76:24]
  wire [2:0] _value_T_3 = deq_ptr_value + 3'h1; // @[Counter.scala 76:24]
  assign ram_class_id_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_class_id_io_deq_bits_MPORT_data = ram_class_id[ram_class_id_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  assign ram_class_id_MPORT_data = io_enq_bits_class_id;
  assign ram_class_id_MPORT_addr = enq_ptr_value;
  assign ram_class_id_MPORT_mask = 1'h1;
  assign ram_class_id_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_host_base_addr_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_host_base_addr_io_deq_bits_MPORT_data = ram_host_base_addr[ram_host_base_addr_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  assign ram_host_base_addr_MPORT_data = io_enq_bits_host_base_addr;
  assign ram_host_base_addr_MPORT_addr = enq_ptr_value;
  assign ram_host_base_addr_MPORT_mask = 1'h1;
  assign ram_host_base_addr_MPORT_en = io_enq_ready & io_enq_valid;
  assign io_enq_ready = ~full; // @[Decoupled.scala 241:19]
  assign io_deq_valid = ~empty; // @[Decoupled.scala 240:19]
  assign io_deq_bits_class_id = ram_class_id_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15]
  assign io_deq_bits_host_base_addr = ram_host_base_addr_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15]
  always @(posedge clock) begin
    if(ram_class_id_MPORT_en & ram_class_id_MPORT_mask) begin
      ram_class_id[ram_class_id_MPORT_addr] <= ram_class_id_MPORT_data; // @[Decoupled.scala 218:16]
    end
    if(ram_host_base_addr_MPORT_en & ram_host_base_addr_MPORT_mask) begin
      ram_host_base_addr[ram_host_base_addr_MPORT_addr] <= ram_host_base_addr_MPORT_data; // @[Decoupled.scala 218:16]
    end
    if (reset) begin // @[Counter.scala 60:40]
      enq_ptr_value <= 3'h0; // @[Counter.scala 60:40]
    end else if (do_enq) begin // @[Decoupled.scala 229:17]
      enq_ptr_value <= _value_T_1; // @[Counter.scala 76:15]
    end
    if (reset) begin // @[Counter.scala 60:40]
      deq_ptr_value <= 3'h0; // @[Counter.scala 60:40]
    end else if (do_deq) begin // @[Decoupled.scala 233:17]
      deq_ptr_value <= _value_T_3; // @[Counter.scala 76:15]
    end
    if (reset) begin // @[Decoupled.scala 221:27]
      maybe_full <= 1'h0; // @[Decoupled.scala 221:27]
    end else if (do_enq != do_deq) begin // @[Decoupled.scala 236:28]
      maybe_full <= do_enq; // @[Decoupled.scala 237:16]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 8; initvar = initvar+1)
    ram_class_id[initvar] = _RAND_0[9:0];
  _RAND_1 = {2{`RANDOM}};
  for (initvar = 0; initvar < 8; initvar = initvar+1)
    ram_host_base_addr[initvar] = _RAND_1[63:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  enq_ptr_value = _RAND_2[2:0];
  _RAND_3 = {1{`RANDOM}};
  deq_ptr_value = _RAND_3[2:0];
  _RAND_4 = {1{`RANDOM}};
  maybe_full = _RAND_4[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module XQueue_2(
  input         clock,
  input         reset,
  output        io_in_ready,
  input         io_in_valid,
  input  [9:0]  io_in_bits_class_id,
  input  [63:0] io_in_bits_host_base_addr,
  input         io_out_ready,
  output        io_out_valid,
  output [9:0]  io_out_bits_class_id,
  output [63:0] io_out_bits_host_base_addr
);
  wire  q_clock; // @[XQueue.scala 85:39]
  wire  q_reset; // @[XQueue.scala 85:39]
  wire  q_io_enq_ready; // @[XQueue.scala 85:39]
  wire  q_io_enq_valid; // @[XQueue.scala 85:39]
  wire [9:0] q_io_enq_bits_class_id; // @[XQueue.scala 85:39]
  wire [63:0] q_io_enq_bits_host_base_addr; // @[XQueue.scala 85:39]
  wire  q_io_deq_ready; // @[XQueue.scala 85:39]
  wire  q_io_deq_valid; // @[XQueue.scala 85:39]
  wire [9:0] q_io_deq_bits_class_id; // @[XQueue.scala 85:39]
  wire [63:0] q_io_deq_bits_host_base_addr; // @[XQueue.scala 85:39]
  Queue_4 q ( // @[XQueue.scala 85:39]
    .clock(q_clock),
    .reset(q_reset),
    .io_enq_ready(q_io_enq_ready),
    .io_enq_valid(q_io_enq_valid),
    .io_enq_bits_class_id(q_io_enq_bits_class_id),
    .io_enq_bits_host_base_addr(q_io_enq_bits_host_base_addr),
    .io_deq_ready(q_io_deq_ready),
    .io_deq_valid(q_io_deq_valid),
    .io_deq_bits_class_id(q_io_deq_bits_class_id),
    .io_deq_bits_host_base_addr(q_io_deq_bits_host_base_addr)
  );
  assign io_in_ready = q_io_enq_ready; // @[XQueue.scala 87:34]
  assign io_out_valid = q_io_deq_valid; // @[XQueue.scala 88:34]
  assign io_out_bits_class_id = q_io_deq_bits_class_id; // @[XQueue.scala 88:34]
  assign io_out_bits_host_base_addr = q_io_deq_bits_host_base_addr; // @[XQueue.scala 88:34]
  assign q_clock = clock;
  assign q_reset = reset;
  assign q_io_enq_valid = io_in_valid; // @[XQueue.scala 87:34]
  assign q_io_enq_bits_class_id = io_in_bits_class_id; // @[XQueue.scala 87:34]
  assign q_io_enq_bits_host_base_addr = io_in_bits_host_base_addr; // @[XQueue.scala 87:34]
  assign q_io_deq_ready = io_out_ready; // @[XQueue.scala 88:34]
endmodule
module Queue_5(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input  [7:0]  io_enq_bits_class_meta_max_field_num,
  input         io_enq_bits_class_meta_field_type_0_is_repeated,
  input  [4:0]  io_enq_bits_class_meta_field_type_0_field_type,
  input  [15:0] io_enq_bits_class_meta_field_type_0_sub_class_id,
  input         io_enq_bits_class_meta_field_type_1_is_repeated,
  input  [4:0]  io_enq_bits_class_meta_field_type_1_field_type,
  input  [15:0] io_enq_bits_class_meta_field_type_1_sub_class_id,
  input         io_enq_bits_class_meta_field_type_2_is_repeated,
  input  [4:0]  io_enq_bits_class_meta_field_type_2_field_type,
  input  [15:0] io_enq_bits_class_meta_field_type_2_sub_class_id,
  input         io_enq_bits_class_meta_field_type_3_is_repeated,
  input  [4:0]  io_enq_bits_class_meta_field_type_3_field_type,
  input  [15:0] io_enq_bits_class_meta_field_type_3_sub_class_id,
  input         io_enq_bits_class_meta_field_type_4_is_repeated,
  input  [4:0]  io_enq_bits_class_meta_field_type_4_field_type,
  input  [15:0] io_enq_bits_class_meta_field_type_4_sub_class_id,
  input         io_enq_bits_class_meta_field_type_5_is_repeated,
  input  [4:0]  io_enq_bits_class_meta_field_type_5_field_type,
  input  [15:0] io_enq_bits_class_meta_field_type_5_sub_class_id,
  input         io_enq_bits_class_meta_field_type_6_is_repeated,
  input  [4:0]  io_enq_bits_class_meta_field_type_6_field_type,
  input  [15:0] io_enq_bits_class_meta_field_type_6_sub_class_id,
  input         io_enq_bits_class_meta_field_type_7_is_repeated,
  input  [4:0]  io_enq_bits_class_meta_field_type_7_field_type,
  input  [15:0] io_enq_bits_class_meta_field_type_7_sub_class_id,
  input         io_enq_bits_class_meta_field_type_8_is_repeated,
  input  [4:0]  io_enq_bits_class_meta_field_type_8_field_type,
  input  [15:0] io_enq_bits_class_meta_field_type_8_sub_class_id,
  input         io_enq_bits_class_meta_field_type_9_is_repeated,
  input  [4:0]  io_enq_bits_class_meta_field_type_9_field_type,
  input  [15:0] io_enq_bits_class_meta_field_type_9_sub_class_id,
  input         io_enq_bits_class_meta_field_type_10_is_repeated,
  input  [4:0]  io_enq_bits_class_meta_field_type_10_field_type,
  input  [15:0] io_enq_bits_class_meta_field_type_10_sub_class_id,
  input         io_enq_bits_class_meta_field_type_11_is_repeated,
  input  [4:0]  io_enq_bits_class_meta_field_type_11_field_type,
  input  [15:0] io_enq_bits_class_meta_field_type_11_sub_class_id,
  input         io_enq_bits_class_meta_field_type_12_is_repeated,
  input  [4:0]  io_enq_bits_class_meta_field_type_12_field_type,
  input  [15:0] io_enq_bits_class_meta_field_type_12_sub_class_id,
  input         io_enq_bits_class_meta_field_type_13_is_repeated,
  input  [4:0]  io_enq_bits_class_meta_field_type_13_field_type,
  input  [15:0] io_enq_bits_class_meta_field_type_13_sub_class_id,
  input         io_enq_bits_class_meta_field_type_14_is_repeated,
  input  [4:0]  io_enq_bits_class_meta_field_type_14_field_type,
  input  [15:0] io_enq_bits_class_meta_field_type_14_sub_class_id,
  input         io_enq_bits_class_meta_field_type_15_is_repeated,
  input  [4:0]  io_enq_bits_class_meta_field_type_15_field_type,
  input  [15:0] io_enq_bits_class_meta_field_type_15_sub_class_id,
  input         io_enq_bits_class_meta_field_type_16_is_repeated,
  input  [4:0]  io_enq_bits_class_meta_field_type_16_field_type,
  input  [15:0] io_enq_bits_class_meta_field_type_16_sub_class_id,
  input         io_enq_bits_class_meta_field_type_17_is_repeated,
  input  [4:0]  io_enq_bits_class_meta_field_type_17_field_type,
  input  [15:0] io_enq_bits_class_meta_field_type_17_sub_class_id,
  input         io_enq_bits_class_meta_field_type_18_is_repeated,
  input  [4:0]  io_enq_bits_class_meta_field_type_18_field_type,
  input  [15:0] io_enq_bits_class_meta_field_type_18_sub_class_id,
  input         io_enq_bits_class_meta_field_type_19_is_repeated,
  input  [4:0]  io_enq_bits_class_meta_field_type_19_field_type,
  input  [15:0] io_enq_bits_class_meta_field_type_19_sub_class_id,
  input         io_enq_bits_class_meta_field_type_20_is_repeated,
  input  [4:0]  io_enq_bits_class_meta_field_type_20_field_type,
  input  [15:0] io_enq_bits_class_meta_field_type_20_sub_class_id,
  input         io_enq_bits_class_meta_field_type_21_is_repeated,
  input  [4:0]  io_enq_bits_class_meta_field_type_21_field_type,
  input  [15:0] io_enq_bits_class_meta_field_type_21_sub_class_id,
  input         io_enq_bits_class_meta_field_type_22_is_repeated,
  input  [4:0]  io_enq_bits_class_meta_field_type_22_field_type,
  input  [15:0] io_enq_bits_class_meta_field_type_22_sub_class_id,
  input         io_enq_bits_class_meta_field_type_23_is_repeated,
  input  [4:0]  io_enq_bits_class_meta_field_type_23_field_type,
  input  [15:0] io_enq_bits_class_meta_field_type_23_sub_class_id,
  input         io_enq_bits_class_meta_field_type_24_is_repeated,
  input  [4:0]  io_enq_bits_class_meta_field_type_24_field_type,
  input  [15:0] io_enq_bits_class_meta_field_type_24_sub_class_id,
  input         io_enq_bits_class_meta_field_type_25_is_repeated,
  input  [4:0]  io_enq_bits_class_meta_field_type_25_field_type,
  input  [15:0] io_enq_bits_class_meta_field_type_25_sub_class_id,
  input         io_enq_bits_class_meta_field_type_26_is_repeated,
  input  [4:0]  io_enq_bits_class_meta_field_type_26_field_type,
  input  [15:0] io_enq_bits_class_meta_field_type_26_sub_class_id,
  input         io_enq_bits_class_meta_field_type_27_is_repeated,
  input  [4:0]  io_enq_bits_class_meta_field_type_27_field_type,
  input  [15:0] io_enq_bits_class_meta_field_type_27_sub_class_id,
  input         io_enq_bits_class_meta_field_type_28_is_repeated,
  input  [4:0]  io_enq_bits_class_meta_field_type_28_field_type,
  input  [15:0] io_enq_bits_class_meta_field_type_28_sub_class_id,
  input         io_enq_bits_class_meta_field_type_29_is_repeated,
  input  [4:0]  io_enq_bits_class_meta_field_type_29_field_type,
  input  [15:0] io_enq_bits_class_meta_field_type_29_sub_class_id,
  input         io_enq_bits_class_meta_field_type_30_is_repeated,
  input  [4:0]  io_enq_bits_class_meta_field_type_30_field_type,
  input  [15:0] io_enq_bits_class_meta_field_type_30_sub_class_id,
  input         io_enq_bits_class_meta_field_type_31_is_repeated,
  input  [4:0]  io_enq_bits_class_meta_field_type_31_field_type,
  input  [15:0] io_enq_bits_class_meta_field_type_31_sub_class_id,
  input         io_enq_bits_class_meta_field_type_32_is_repeated,
  input  [4:0]  io_enq_bits_class_meta_field_type_32_field_type,
  input  [15:0] io_enq_bits_class_meta_field_type_32_sub_class_id,
  input         io_deq_ready,
  output        io_deq_valid,
  output [7:0]  io_deq_bits_class_meta_max_field_num,
  output        io_deq_bits_class_meta_field_type_0_is_repeated,
  output [4:0]  io_deq_bits_class_meta_field_type_0_field_type,
  output [15:0] io_deq_bits_class_meta_field_type_0_sub_class_id,
  output        io_deq_bits_class_meta_field_type_1_is_repeated,
  output [4:0]  io_deq_bits_class_meta_field_type_1_field_type,
  output [15:0] io_deq_bits_class_meta_field_type_1_sub_class_id,
  output        io_deq_bits_class_meta_field_type_2_is_repeated,
  output [4:0]  io_deq_bits_class_meta_field_type_2_field_type,
  output [15:0] io_deq_bits_class_meta_field_type_2_sub_class_id,
  output        io_deq_bits_class_meta_field_type_3_is_repeated,
  output [4:0]  io_deq_bits_class_meta_field_type_3_field_type,
  output [15:0] io_deq_bits_class_meta_field_type_3_sub_class_id,
  output        io_deq_bits_class_meta_field_type_4_is_repeated,
  output [4:0]  io_deq_bits_class_meta_field_type_4_field_type,
  output [15:0] io_deq_bits_class_meta_field_type_4_sub_class_id,
  output        io_deq_bits_class_meta_field_type_5_is_repeated,
  output [4:0]  io_deq_bits_class_meta_field_type_5_field_type,
  output [15:0] io_deq_bits_class_meta_field_type_5_sub_class_id,
  output        io_deq_bits_class_meta_field_type_6_is_repeated,
  output [4:0]  io_deq_bits_class_meta_field_type_6_field_type,
  output [15:0] io_deq_bits_class_meta_field_type_6_sub_class_id,
  output        io_deq_bits_class_meta_field_type_7_is_repeated,
  output [4:0]  io_deq_bits_class_meta_field_type_7_field_type,
  output [15:0] io_deq_bits_class_meta_field_type_7_sub_class_id,
  output        io_deq_bits_class_meta_field_type_8_is_repeated,
  output [4:0]  io_deq_bits_class_meta_field_type_8_field_type,
  output [15:0] io_deq_bits_class_meta_field_type_8_sub_class_id,
  output        io_deq_bits_class_meta_field_type_9_is_repeated,
  output [4:0]  io_deq_bits_class_meta_field_type_9_field_type,
  output [15:0] io_deq_bits_class_meta_field_type_9_sub_class_id,
  output        io_deq_bits_class_meta_field_type_10_is_repeated,
  output [4:0]  io_deq_bits_class_meta_field_type_10_field_type,
  output [15:0] io_deq_bits_class_meta_field_type_10_sub_class_id,
  output        io_deq_bits_class_meta_field_type_11_is_repeated,
  output [4:0]  io_deq_bits_class_meta_field_type_11_field_type,
  output [15:0] io_deq_bits_class_meta_field_type_11_sub_class_id,
  output        io_deq_bits_class_meta_field_type_12_is_repeated,
  output [4:0]  io_deq_bits_class_meta_field_type_12_field_type,
  output [15:0] io_deq_bits_class_meta_field_type_12_sub_class_id,
  output        io_deq_bits_class_meta_field_type_13_is_repeated,
  output [4:0]  io_deq_bits_class_meta_field_type_13_field_type,
  output [15:0] io_deq_bits_class_meta_field_type_13_sub_class_id,
  output        io_deq_bits_class_meta_field_type_14_is_repeated,
  output [4:0]  io_deq_bits_class_meta_field_type_14_field_type,
  output [15:0] io_deq_bits_class_meta_field_type_14_sub_class_id,
  output        io_deq_bits_class_meta_field_type_15_is_repeated,
  output [4:0]  io_deq_bits_class_meta_field_type_15_field_type,
  output [15:0] io_deq_bits_class_meta_field_type_15_sub_class_id,
  output        io_deq_bits_class_meta_field_type_16_is_repeated,
  output [4:0]  io_deq_bits_class_meta_field_type_16_field_type,
  output [15:0] io_deq_bits_class_meta_field_type_16_sub_class_id,
  output        io_deq_bits_class_meta_field_type_17_is_repeated,
  output [4:0]  io_deq_bits_class_meta_field_type_17_field_type,
  output [15:0] io_deq_bits_class_meta_field_type_17_sub_class_id,
  output        io_deq_bits_class_meta_field_type_18_is_repeated,
  output [4:0]  io_deq_bits_class_meta_field_type_18_field_type,
  output [15:0] io_deq_bits_class_meta_field_type_18_sub_class_id,
  output        io_deq_bits_class_meta_field_type_19_is_repeated,
  output [4:0]  io_deq_bits_class_meta_field_type_19_field_type,
  output [15:0] io_deq_bits_class_meta_field_type_19_sub_class_id,
  output        io_deq_bits_class_meta_field_type_20_is_repeated,
  output [4:0]  io_deq_bits_class_meta_field_type_20_field_type,
  output [15:0] io_deq_bits_class_meta_field_type_20_sub_class_id,
  output        io_deq_bits_class_meta_field_type_21_is_repeated,
  output [4:0]  io_deq_bits_class_meta_field_type_21_field_type,
  output [15:0] io_deq_bits_class_meta_field_type_21_sub_class_id,
  output        io_deq_bits_class_meta_field_type_22_is_repeated,
  output [4:0]  io_deq_bits_class_meta_field_type_22_field_type,
  output [15:0] io_deq_bits_class_meta_field_type_22_sub_class_id,
  output        io_deq_bits_class_meta_field_type_23_is_repeated,
  output [4:0]  io_deq_bits_class_meta_field_type_23_field_type,
  output [15:0] io_deq_bits_class_meta_field_type_23_sub_class_id,
  output        io_deq_bits_class_meta_field_type_24_is_repeated,
  output [4:0]  io_deq_bits_class_meta_field_type_24_field_type,
  output [15:0] io_deq_bits_class_meta_field_type_24_sub_class_id,
  output        io_deq_bits_class_meta_field_type_25_is_repeated,
  output [4:0]  io_deq_bits_class_meta_field_type_25_field_type,
  output [15:0] io_deq_bits_class_meta_field_type_25_sub_class_id,
  output        io_deq_bits_class_meta_field_type_26_is_repeated,
  output [4:0]  io_deq_bits_class_meta_field_type_26_field_type,
  output [15:0] io_deq_bits_class_meta_field_type_26_sub_class_id,
  output        io_deq_bits_class_meta_field_type_27_is_repeated,
  output [4:0]  io_deq_bits_class_meta_field_type_27_field_type,
  output [15:0] io_deq_bits_class_meta_field_type_27_sub_class_id,
  output        io_deq_bits_class_meta_field_type_28_is_repeated,
  output [4:0]  io_deq_bits_class_meta_field_type_28_field_type,
  output [15:0] io_deq_bits_class_meta_field_type_28_sub_class_id,
  output        io_deq_bits_class_meta_field_type_29_is_repeated,
  output [4:0]  io_deq_bits_class_meta_field_type_29_field_type,
  output [15:0] io_deq_bits_class_meta_field_type_29_sub_class_id,
  output        io_deq_bits_class_meta_field_type_30_is_repeated,
  output [4:0]  io_deq_bits_class_meta_field_type_30_field_type,
  output [15:0] io_deq_bits_class_meta_field_type_30_sub_class_id,
  output        io_deq_bits_class_meta_field_type_31_is_repeated,
  output [4:0]  io_deq_bits_class_meta_field_type_31_field_type,
  output [15:0] io_deq_bits_class_meta_field_type_31_sub_class_id,
  output        io_deq_bits_class_meta_field_type_32_is_repeated,
  output [4:0]  io_deq_bits_class_meta_field_type_32_field_type,
  output [15:0] io_deq_bits_class_meta_field_type_32_sub_class_id
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
`endif // RANDOMIZE_REG_INIT
  reg [7:0] ram_class_meta_max_field_num [0:7]; // @[Decoupled.scala 218:16]
  wire [7:0] ram_class_meta_max_field_num_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16]
  wire [2:0] ram_class_meta_max_field_num_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16]
  wire [7:0] ram_class_meta_max_field_num_MPORT_data; // @[Decoupled.scala 218:16]
  wire [2:0] ram_class_meta_max_field_num_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_class_meta_max_field_num_MPORT_mask; // @[Decoupled.scala 218:16]
  wire  ram_class_meta_max_field_num_MPORT_en; // @[Decoupled.scala 218:16]
  reg  ram_class_meta_field_type_0_is_repeated [0:7]; // @[Decoupled.scala 218:16]
  wire  ram_class_meta_field_type_0_is_repeated_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16]
  wire [2:0] ram_class_meta_field_type_0_is_repeated_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_class_meta_field_type_0_is_repeated_MPORT_data; // @[Decoupled.scala 218:16]
  wire [2:0] ram_class_meta_field_type_0_is_repeated_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_class_meta_field_type_0_is_repeated_MPORT_mask; // @[Decoupled.scala 218:16]
  wire  ram_class_meta_field_type_0_is_repeated_MPORT_en; // @[Decoupled.scala 218:16]
  reg [4:0] ram_class_meta_field_type_0_field_type [0:7]; // @[Decoupled.scala 218:16]
  wire [4:0] ram_class_meta_field_type_0_field_type_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16]
  wire [2:0] ram_class_meta_field_type_0_field_type_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16]
  wire [4:0] ram_class_meta_field_type_0_field_type_MPORT_data; // @[Decoupled.scala 218:16]
  wire [2:0] ram_class_meta_field_type_0_field_type_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_class_meta_field_type_0_field_type_MPORT_mask; // @[Decoupled.scala 218:16]
  wire  ram_class_meta_field_type_0_field_type_MPORT_en; // @[Decoupled.scala 218:16]
  reg [15:0] ram_class_meta_field_type_0_sub_class_id [0:7]; // @[Decoupled.scala 218:16]
  wire [15:0] ram_class_meta_field_type_0_sub_class_id_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16]
  wire [2:0] ram_class_meta_field_type_0_sub_class_id_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16]
  wire [15:0] ram_class_meta_field_type_0_sub_class_id_MPORT_data; // @[Decoupled.scala 218:16]
  wire [2:0] ram_class_meta_field_type_0_sub_class_id_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_class_meta_field_type_0_sub_class_id_MPORT_mask; // @[Decoupled.scala 218:16]
  wire  ram_class_meta_field_type_0_sub_class_id_MPORT_en; // @[Decoupled.scala 218:16]
  reg  ram_class_meta_field_type_1_is_repeated [0:7]; // @[Decoupled.scala 218:16]
  wire  ram_class_meta_field_type_1_is_repeated_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16]
  wire [2:0] ram_class_meta_field_type_1_is_repeated_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_class_meta_field_type_1_is_repeated_MPORT_data; // @[Decoupled.scala 218:16]
  wire [2:0] ram_class_meta_field_type_1_is_repeated_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_class_meta_field_type_1_is_repeated_MPORT_mask; // @[Decoupled.scala 218:16]
  wire  ram_class_meta_field_type_1_is_repeated_MPORT_en; // @[Decoupled.scala 218:16]
  reg [4:0] ram_class_meta_field_type_1_field_type [0:7]; // @[Decoupled.scala 218:16]
  wire [4:0] ram_class_meta_field_type_1_field_type_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16]
  wire [2:0] ram_class_meta_field_type_1_field_type_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16]
  wire [4:0] ram_class_meta_field_type_1_field_type_MPORT_data; // @[Decoupled.scala 218:16]
  wire [2:0] ram_class_meta_field_type_1_field_type_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_class_meta_field_type_1_field_type_MPORT_mask; // @[Decoupled.scala 218:16]
  wire  ram_class_meta_field_type_1_field_type_MPORT_en; // @[Decoupled.scala 218:16]
  reg [15:0] ram_class_meta_field_type_1_sub_class_id [0:7]; // @[Decoupled.scala 218:16]
  wire [15:0] ram_class_meta_field_type_1_sub_class_id_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16]
  wire [2:0] ram_class_meta_field_type_1_sub_class_id_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16]
  wire [15:0] ram_class_meta_field_type_1_sub_class_id_MPORT_data; // @[Decoupled.scala 218:16]
  wire [2:0] ram_class_meta_field_type_1_sub_class_id_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_class_meta_field_type_1_sub_class_id_MPORT_mask; // @[Decoupled.scala 218:16]
  wire  ram_class_meta_field_type_1_sub_class_id_MPORT_en; // @[Decoupled.scala 218:16]
  reg  ram_class_meta_field_type_2_is_repeated [0:7]; // @[Decoupled.scala 218:16]
  wire  ram_class_meta_field_type_2_is_repeated_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16]
  wire [2:0] ram_class_meta_field_type_2_is_repeated_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_class_meta_field_type_2_is_repeated_MPORT_data; // @[Decoupled.scala 218:16]
  wire [2:0] ram_class_meta_field_type_2_is_repeated_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_class_meta_field_type_2_is_repeated_MPORT_mask; // @[Decoupled.scala 218:16]
  wire  ram_class_meta_field_type_2_is_repeated_MPORT_en; // @[Decoupled.scala 218:16]
  reg [4:0] ram_class_meta_field_type_2_field_type [0:7]; // @[Decoupled.scala 218:16]
  wire [4:0] ram_class_meta_field_type_2_field_type_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16]
  wire [2:0] ram_class_meta_field_type_2_field_type_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16]
  wire [4:0] ram_class_meta_field_type_2_field_type_MPORT_data; // @[Decoupled.scala 218:16]
  wire [2:0] ram_class_meta_field_type_2_field_type_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_class_meta_field_type_2_field_type_MPORT_mask; // @[Decoupled.scala 218:16]
  wire  ram_class_meta_field_type_2_field_type_MPORT_en; // @[Decoupled.scala 218:16]
  reg [15:0] ram_class_meta_field_type_2_sub_class_id [0:7]; // @[Decoupled.scala 218:16]
  wire [15:0] ram_class_meta_field_type_2_sub_class_id_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16]
  wire [2:0] ram_class_meta_field_type_2_sub_class_id_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16]
  wire [15:0] ram_class_meta_field_type_2_sub_class_id_MPORT_data; // @[Decoupled.scala 218:16]
  wire [2:0] ram_class_meta_field_type_2_sub_class_id_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_class_meta_field_type_2_sub_class_id_MPORT_mask; // @[Decoupled.scala 218:16]
  wire  ram_class_meta_field_type_2_sub_class_id_MPORT_en; // @[Decoupled.scala 218:16]
  reg  ram_class_meta_field_type_3_is_repeated [0:7]; // @[Decoupled.scala 218:16]
  wire  ram_class_meta_field_type_3_is_repeated_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16]
  wire [2:0] ram_class_meta_field_type_3_is_repeated_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_class_meta_field_type_3_is_repeated_MPORT_data; // @[Decoupled.scala 218:16]
  wire [2:0] ram_class_meta_field_type_3_is_repeated_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_class_meta_field_type_3_is_repeated_MPORT_mask; // @[Decoupled.scala 218:16]
  wire  ram_class_meta_field_type_3_is_repeated_MPORT_en; // @[Decoupled.scala 218:16]
  reg [4:0] ram_class_meta_field_type_3_field_type [0:7]; // @[Decoupled.scala 218:16]
  wire [4:0] ram_class_meta_field_type_3_field_type_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16]
  wire [2:0] ram_class_meta_field_type_3_field_type_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16]
  wire [4:0] ram_class_meta_field_type_3_field_type_MPORT_data; // @[Decoupled.scala 218:16]
  wire [2:0] ram_class_meta_field_type_3_field_type_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_class_meta_field_type_3_field_type_MPORT_mask; // @[Decoupled.scala 218:16]
  wire  ram_class_meta_field_type_3_field_type_MPORT_en; // @[Decoupled.scala 218:16]
  reg [15:0] ram_class_meta_field_type_3_sub_class_id [0:7]; // @[Decoupled.scala 218:16]
  wire [15:0] ram_class_meta_field_type_3_sub_class_id_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16]
  wire [2:0] ram_class_meta_field_type_3_sub_class_id_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16]
  wire [15:0] ram_class_meta_field_type_3_sub_class_id_MPORT_data; // @[Decoupled.scala 218:16]
  wire [2:0] ram_class_meta_field_type_3_sub_class_id_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_class_meta_field_type_3_sub_class_id_MPORT_mask; // @[Decoupled.scala 218:16]
  wire  ram_class_meta_field_type_3_sub_class_id_MPORT_en; // @[Decoupled.scala 218:16]
  reg  ram_class_meta_field_type_4_is_repeated [0:7]; // @[Decoupled.scala 218:16]
  wire  ram_class_meta_field_type_4_is_repeated_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16]
  wire [2:0] ram_class_meta_field_type_4_is_repeated_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_class_meta_field_type_4_is_repeated_MPORT_data; // @[Decoupled.scala 218:16]
  wire [2:0] ram_class_meta_field_type_4_is_repeated_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_class_meta_field_type_4_is_repeated_MPORT_mask; // @[Decoupled.scala 218:16]
  wire  ram_class_meta_field_type_4_is_repeated_MPORT_en; // @[Decoupled.scala 218:16]
  reg [4:0] ram_class_meta_field_type_4_field_type [0:7]; // @[Decoupled.scala 218:16]
  wire [4:0] ram_class_meta_field_type_4_field_type_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16]
  wire [2:0] ram_class_meta_field_type_4_field_type_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16]
  wire [4:0] ram_class_meta_field_type_4_field_type_MPORT_data; // @[Decoupled.scala 218:16]
  wire [2:0] ram_class_meta_field_type_4_field_type_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_class_meta_field_type_4_field_type_MPORT_mask; // @[Decoupled.scala 218:16]
  wire  ram_class_meta_field_type_4_field_type_MPORT_en; // @[Decoupled.scala 218:16]
  reg [15:0] ram_class_meta_field_type_4_sub_class_id [0:7]; // @[Decoupled.scala 218:16]
  wire [15:0] ram_class_meta_field_type_4_sub_class_id_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16]
  wire [2:0] ram_class_meta_field_type_4_sub_class_id_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16]
  wire [15:0] ram_class_meta_field_type_4_sub_class_id_MPORT_data; // @[Decoupled.scala 218:16]
  wire [2:0] ram_class_meta_field_type_4_sub_class_id_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_class_meta_field_type_4_sub_class_id_MPORT_mask; // @[Decoupled.scala 218:16]
  wire  ram_class_meta_field_type_4_sub_class_id_MPORT_en; // @[Decoupled.scala 218:16]
  reg  ram_class_meta_field_type_5_is_repeated [0:7]; // @[Decoupled.scala 218:16]
  wire  ram_class_meta_field_type_5_is_repeated_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16]
  wire [2:0] ram_class_meta_field_type_5_is_repeated_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_class_meta_field_type_5_is_repeated_MPORT_data; // @[Decoupled.scala 218:16]
  wire [2:0] ram_class_meta_field_type_5_is_repeated_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_class_meta_field_type_5_is_repeated_MPORT_mask; // @[Decoupled.scala 218:16]
  wire  ram_class_meta_field_type_5_is_repeated_MPORT_en; // @[Decoupled.scala 218:16]
  reg [4:0] ram_class_meta_field_type_5_field_type [0:7]; // @[Decoupled.scala 218:16]
  wire [4:0] ram_class_meta_field_type_5_field_type_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16]
  wire [2:0] ram_class_meta_field_type_5_field_type_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16]
  wire [4:0] ram_class_meta_field_type_5_field_type_MPORT_data; // @[Decoupled.scala 218:16]
  wire [2:0] ram_class_meta_field_type_5_field_type_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_class_meta_field_type_5_field_type_MPORT_mask; // @[Decoupled.scala 218:16]
  wire  ram_class_meta_field_type_5_field_type_MPORT_en; // @[Decoupled.scala 218:16]
  reg [15:0] ram_class_meta_field_type_5_sub_class_id [0:7]; // @[Decoupled.scala 218:16]
  wire [15:0] ram_class_meta_field_type_5_sub_class_id_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16]
  wire [2:0] ram_class_meta_field_type_5_sub_class_id_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16]
  wire [15:0] ram_class_meta_field_type_5_sub_class_id_MPORT_data; // @[Decoupled.scala 218:16]
  wire [2:0] ram_class_meta_field_type_5_sub_class_id_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_class_meta_field_type_5_sub_class_id_MPORT_mask; // @[Decoupled.scala 218:16]
  wire  ram_class_meta_field_type_5_sub_class_id_MPORT_en; // @[Decoupled.scala 218:16]
  reg  ram_class_meta_field_type_6_is_repeated [0:7]; // @[Decoupled.scala 218:16]
  wire  ram_class_meta_field_type_6_is_repeated_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16]
  wire [2:0] ram_class_meta_field_type_6_is_repeated_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_class_meta_field_type_6_is_repeated_MPORT_data; // @[Decoupled.scala 218:16]
  wire [2:0] ram_class_meta_field_type_6_is_repeated_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_class_meta_field_type_6_is_repeated_MPORT_mask; // @[Decoupled.scala 218:16]
  wire  ram_class_meta_field_type_6_is_repeated_MPORT_en; // @[Decoupled.scala 218:16]
  reg [4:0] ram_class_meta_field_type_6_field_type [0:7]; // @[Decoupled.scala 218:16]
  wire [4:0] ram_class_meta_field_type_6_field_type_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16]
  wire [2:0] ram_class_meta_field_type_6_field_type_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16]
  wire [4:0] ram_class_meta_field_type_6_field_type_MPORT_data; // @[Decoupled.scala 218:16]
  wire [2:0] ram_class_meta_field_type_6_field_type_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_class_meta_field_type_6_field_type_MPORT_mask; // @[Decoupled.scala 218:16]
  wire  ram_class_meta_field_type_6_field_type_MPORT_en; // @[Decoupled.scala 218:16]
  reg [15:0] ram_class_meta_field_type_6_sub_class_id [0:7]; // @[Decoupled.scala 218:16]
  wire [15:0] ram_class_meta_field_type_6_sub_class_id_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16]
  wire [2:0] ram_class_meta_field_type_6_sub_class_id_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16]
  wire [15:0] ram_class_meta_field_type_6_sub_class_id_MPORT_data; // @[Decoupled.scala 218:16]
  wire [2:0] ram_class_meta_field_type_6_sub_class_id_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_class_meta_field_type_6_sub_class_id_MPORT_mask; // @[Decoupled.scala 218:16]
  wire  ram_class_meta_field_type_6_sub_class_id_MPORT_en; // @[Decoupled.scala 218:16]
  reg  ram_class_meta_field_type_7_is_repeated [0:7]; // @[Decoupled.scala 218:16]
  wire  ram_class_meta_field_type_7_is_repeated_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16]
  wire [2:0] ram_class_meta_field_type_7_is_repeated_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_class_meta_field_type_7_is_repeated_MPORT_data; // @[Decoupled.scala 218:16]
  wire [2:0] ram_class_meta_field_type_7_is_repeated_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_class_meta_field_type_7_is_repeated_MPORT_mask; // @[Decoupled.scala 218:16]
  wire  ram_class_meta_field_type_7_is_repeated_MPORT_en; // @[Decoupled.scala 218:16]
  reg [4:0] ram_class_meta_field_type_7_field_type [0:7]; // @[Decoupled.scala 218:16]
  wire [4:0] ram_class_meta_field_type_7_field_type_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16]
  wire [2:0] ram_class_meta_field_type_7_field_type_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16]
  wire [4:0] ram_class_meta_field_type_7_field_type_MPORT_data; // @[Decoupled.scala 218:16]
  wire [2:0] ram_class_meta_field_type_7_field_type_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_class_meta_field_type_7_field_type_MPORT_mask; // @[Decoupled.scala 218:16]
  wire  ram_class_meta_field_type_7_field_type_MPORT_en; // @[Decoupled.scala 218:16]
  reg [15:0] ram_class_meta_field_type_7_sub_class_id [0:7]; // @[Decoupled.scala 218:16]
  wire [15:0] ram_class_meta_field_type_7_sub_class_id_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16]
  wire [2:0] ram_class_meta_field_type_7_sub_class_id_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16]
  wire [15:0] ram_class_meta_field_type_7_sub_class_id_MPORT_data; // @[Decoupled.scala 218:16]
  wire [2:0] ram_class_meta_field_type_7_sub_class_id_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_class_meta_field_type_7_sub_class_id_MPORT_mask; // @[Decoupled.scala 218:16]
  wire  ram_class_meta_field_type_7_sub_class_id_MPORT_en; // @[Decoupled.scala 218:16]
  reg  ram_class_meta_field_type_8_is_repeated [0:7]; // @[Decoupled.scala 218:16]
  wire  ram_class_meta_field_type_8_is_repeated_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16]
  wire [2:0] ram_class_meta_field_type_8_is_repeated_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_class_meta_field_type_8_is_repeated_MPORT_data; // @[Decoupled.scala 218:16]
  wire [2:0] ram_class_meta_field_type_8_is_repeated_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_class_meta_field_type_8_is_repeated_MPORT_mask; // @[Decoupled.scala 218:16]
  wire  ram_class_meta_field_type_8_is_repeated_MPORT_en; // @[Decoupled.scala 218:16]
  reg [4:0] ram_class_meta_field_type_8_field_type [0:7]; // @[Decoupled.scala 218:16]
  wire [4:0] ram_class_meta_field_type_8_field_type_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16]
  wire [2:0] ram_class_meta_field_type_8_field_type_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16]
  wire [4:0] ram_class_meta_field_type_8_field_type_MPORT_data; // @[Decoupled.scala 218:16]
  wire [2:0] ram_class_meta_field_type_8_field_type_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_class_meta_field_type_8_field_type_MPORT_mask; // @[Decoupled.scala 218:16]
  wire  ram_class_meta_field_type_8_field_type_MPORT_en; // @[Decoupled.scala 218:16]
  reg [15:0] ram_class_meta_field_type_8_sub_class_id [0:7]; // @[Decoupled.scala 218:16]
  wire [15:0] ram_class_meta_field_type_8_sub_class_id_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16]
  wire [2:0] ram_class_meta_field_type_8_sub_class_id_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16]
  wire [15:0] ram_class_meta_field_type_8_sub_class_id_MPORT_data; // @[Decoupled.scala 218:16]
  wire [2:0] ram_class_meta_field_type_8_sub_class_id_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_class_meta_field_type_8_sub_class_id_MPORT_mask; // @[Decoupled.scala 218:16]
  wire  ram_class_meta_field_type_8_sub_class_id_MPORT_en; // @[Decoupled.scala 218:16]
  reg  ram_class_meta_field_type_9_is_repeated [0:7]; // @[Decoupled.scala 218:16]
  wire  ram_class_meta_field_type_9_is_repeated_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16]
  wire [2:0] ram_class_meta_field_type_9_is_repeated_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_class_meta_field_type_9_is_repeated_MPORT_data; // @[Decoupled.scala 218:16]
  wire [2:0] ram_class_meta_field_type_9_is_repeated_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_class_meta_field_type_9_is_repeated_MPORT_mask; // @[Decoupled.scala 218:16]
  wire  ram_class_meta_field_type_9_is_repeated_MPORT_en; // @[Decoupled.scala 218:16]
  reg [4:0] ram_class_meta_field_type_9_field_type [0:7]; // @[Decoupled.scala 218:16]
  wire [4:0] ram_class_meta_field_type_9_field_type_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16]
  wire [2:0] ram_class_meta_field_type_9_field_type_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16]
  wire [4:0] ram_class_meta_field_type_9_field_type_MPORT_data; // @[Decoupled.scala 218:16]
  wire [2:0] ram_class_meta_field_type_9_field_type_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_class_meta_field_type_9_field_type_MPORT_mask; // @[Decoupled.scala 218:16]
  wire  ram_class_meta_field_type_9_field_type_MPORT_en; // @[Decoupled.scala 218:16]
  reg [15:0] ram_class_meta_field_type_9_sub_class_id [0:7]; // @[Decoupled.scala 218:16]
  wire [15:0] ram_class_meta_field_type_9_sub_class_id_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16]
  wire [2:0] ram_class_meta_field_type_9_sub_class_id_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16]
  wire [15:0] ram_class_meta_field_type_9_sub_class_id_MPORT_data; // @[Decoupled.scala 218:16]
  wire [2:0] ram_class_meta_field_type_9_sub_class_id_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_class_meta_field_type_9_sub_class_id_MPORT_mask; // @[Decoupled.scala 218:16]
  wire  ram_class_meta_field_type_9_sub_class_id_MPORT_en; // @[Decoupled.scala 218:16]
  reg  ram_class_meta_field_type_10_is_repeated [0:7]; // @[Decoupled.scala 218:16]
  wire  ram_class_meta_field_type_10_is_repeated_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16]
  wire [2:0] ram_class_meta_field_type_10_is_repeated_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_class_meta_field_type_10_is_repeated_MPORT_data; // @[Decoupled.scala 218:16]
  wire [2:0] ram_class_meta_field_type_10_is_repeated_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_class_meta_field_type_10_is_repeated_MPORT_mask; // @[Decoupled.scala 218:16]
  wire  ram_class_meta_field_type_10_is_repeated_MPORT_en; // @[Decoupled.scala 218:16]
  reg [4:0] ram_class_meta_field_type_10_field_type [0:7]; // @[Decoupled.scala 218:16]
  wire [4:0] ram_class_meta_field_type_10_field_type_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16]
  wire [2:0] ram_class_meta_field_type_10_field_type_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16]
  wire [4:0] ram_class_meta_field_type_10_field_type_MPORT_data; // @[Decoupled.scala 218:16]
  wire [2:0] ram_class_meta_field_type_10_field_type_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_class_meta_field_type_10_field_type_MPORT_mask; // @[Decoupled.scala 218:16]
  wire  ram_class_meta_field_type_10_field_type_MPORT_en; // @[Decoupled.scala 218:16]
  reg [15:0] ram_class_meta_field_type_10_sub_class_id [0:7]; // @[Decoupled.scala 218:16]
  wire [15:0] ram_class_meta_field_type_10_sub_class_id_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16]
  wire [2:0] ram_class_meta_field_type_10_sub_class_id_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16]
  wire [15:0] ram_class_meta_field_type_10_sub_class_id_MPORT_data; // @[Decoupled.scala 218:16]
  wire [2:0] ram_class_meta_field_type_10_sub_class_id_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_class_meta_field_type_10_sub_class_id_MPORT_mask; // @[Decoupled.scala 218:16]
  wire  ram_class_meta_field_type_10_sub_class_id_MPORT_en; // @[Decoupled.scala 218:16]
  reg  ram_class_meta_field_type_11_is_repeated [0:7]; // @[Decoupled.scala 218:16]
  wire  ram_class_meta_field_type_11_is_repeated_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16]
  wire [2:0] ram_class_meta_field_type_11_is_repeated_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_class_meta_field_type_11_is_repeated_MPORT_data; // @[Decoupled.scala 218:16]
  wire [2:0] ram_class_meta_field_type_11_is_repeated_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_class_meta_field_type_11_is_repeated_MPORT_mask; // @[Decoupled.scala 218:16]
  wire  ram_class_meta_field_type_11_is_repeated_MPORT_en; // @[Decoupled.scala 218:16]
  reg [4:0] ram_class_meta_field_type_11_field_type [0:7]; // @[Decoupled.scala 218:16]
  wire [4:0] ram_class_meta_field_type_11_field_type_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16]
  wire [2:0] ram_class_meta_field_type_11_field_type_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16]
  wire [4:0] ram_class_meta_field_type_11_field_type_MPORT_data; // @[Decoupled.scala 218:16]
  wire [2:0] ram_class_meta_field_type_11_field_type_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_class_meta_field_type_11_field_type_MPORT_mask; // @[Decoupled.scala 218:16]
  wire  ram_class_meta_field_type_11_field_type_MPORT_en; // @[Decoupled.scala 218:16]
  reg [15:0] ram_class_meta_field_type_11_sub_class_id [0:7]; // @[Decoupled.scala 218:16]
  wire [15:0] ram_class_meta_field_type_11_sub_class_id_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16]
  wire [2:0] ram_class_meta_field_type_11_sub_class_id_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16]
  wire [15:0] ram_class_meta_field_type_11_sub_class_id_MPORT_data; // @[Decoupled.scala 218:16]
  wire [2:0] ram_class_meta_field_type_11_sub_class_id_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_class_meta_field_type_11_sub_class_id_MPORT_mask; // @[Decoupled.scala 218:16]
  wire  ram_class_meta_field_type_11_sub_class_id_MPORT_en; // @[Decoupled.scala 218:16]
  reg  ram_class_meta_field_type_12_is_repeated [0:7]; // @[Decoupled.scala 218:16]
  wire  ram_class_meta_field_type_12_is_repeated_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16]
  wire [2:0] ram_class_meta_field_type_12_is_repeated_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_class_meta_field_type_12_is_repeated_MPORT_data; // @[Decoupled.scala 218:16]
  wire [2:0] ram_class_meta_field_type_12_is_repeated_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_class_meta_field_type_12_is_repeated_MPORT_mask; // @[Decoupled.scala 218:16]
  wire  ram_class_meta_field_type_12_is_repeated_MPORT_en; // @[Decoupled.scala 218:16]
  reg [4:0] ram_class_meta_field_type_12_field_type [0:7]; // @[Decoupled.scala 218:16]
  wire [4:0] ram_class_meta_field_type_12_field_type_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16]
  wire [2:0] ram_class_meta_field_type_12_field_type_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16]
  wire [4:0] ram_class_meta_field_type_12_field_type_MPORT_data; // @[Decoupled.scala 218:16]
  wire [2:0] ram_class_meta_field_type_12_field_type_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_class_meta_field_type_12_field_type_MPORT_mask; // @[Decoupled.scala 218:16]
  wire  ram_class_meta_field_type_12_field_type_MPORT_en; // @[Decoupled.scala 218:16]
  reg [15:0] ram_class_meta_field_type_12_sub_class_id [0:7]; // @[Decoupled.scala 218:16]
  wire [15:0] ram_class_meta_field_type_12_sub_class_id_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16]
  wire [2:0] ram_class_meta_field_type_12_sub_class_id_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16]
  wire [15:0] ram_class_meta_field_type_12_sub_class_id_MPORT_data; // @[Decoupled.scala 218:16]
  wire [2:0] ram_class_meta_field_type_12_sub_class_id_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_class_meta_field_type_12_sub_class_id_MPORT_mask; // @[Decoupled.scala 218:16]
  wire  ram_class_meta_field_type_12_sub_class_id_MPORT_en; // @[Decoupled.scala 218:16]
  reg  ram_class_meta_field_type_13_is_repeated [0:7]; // @[Decoupled.scala 218:16]
  wire  ram_class_meta_field_type_13_is_repeated_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16]
  wire [2:0] ram_class_meta_field_type_13_is_repeated_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_class_meta_field_type_13_is_repeated_MPORT_data; // @[Decoupled.scala 218:16]
  wire [2:0] ram_class_meta_field_type_13_is_repeated_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_class_meta_field_type_13_is_repeated_MPORT_mask; // @[Decoupled.scala 218:16]
  wire  ram_class_meta_field_type_13_is_repeated_MPORT_en; // @[Decoupled.scala 218:16]
  reg [4:0] ram_class_meta_field_type_13_field_type [0:7]; // @[Decoupled.scala 218:16]
  wire [4:0] ram_class_meta_field_type_13_field_type_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16]
  wire [2:0] ram_class_meta_field_type_13_field_type_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16]
  wire [4:0] ram_class_meta_field_type_13_field_type_MPORT_data; // @[Decoupled.scala 218:16]
  wire [2:0] ram_class_meta_field_type_13_field_type_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_class_meta_field_type_13_field_type_MPORT_mask; // @[Decoupled.scala 218:16]
  wire  ram_class_meta_field_type_13_field_type_MPORT_en; // @[Decoupled.scala 218:16]
  reg [15:0] ram_class_meta_field_type_13_sub_class_id [0:7]; // @[Decoupled.scala 218:16]
  wire [15:0] ram_class_meta_field_type_13_sub_class_id_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16]
  wire [2:0] ram_class_meta_field_type_13_sub_class_id_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16]
  wire [15:0] ram_class_meta_field_type_13_sub_class_id_MPORT_data; // @[Decoupled.scala 218:16]
  wire [2:0] ram_class_meta_field_type_13_sub_class_id_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_class_meta_field_type_13_sub_class_id_MPORT_mask; // @[Decoupled.scala 218:16]
  wire  ram_class_meta_field_type_13_sub_class_id_MPORT_en; // @[Decoupled.scala 218:16]
  reg  ram_class_meta_field_type_14_is_repeated [0:7]; // @[Decoupled.scala 218:16]
  wire  ram_class_meta_field_type_14_is_repeated_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16]
  wire [2:0] ram_class_meta_field_type_14_is_repeated_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_class_meta_field_type_14_is_repeated_MPORT_data; // @[Decoupled.scala 218:16]
  wire [2:0] ram_class_meta_field_type_14_is_repeated_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_class_meta_field_type_14_is_repeated_MPORT_mask; // @[Decoupled.scala 218:16]
  wire  ram_class_meta_field_type_14_is_repeated_MPORT_en; // @[Decoupled.scala 218:16]
  reg [4:0] ram_class_meta_field_type_14_field_type [0:7]; // @[Decoupled.scala 218:16]
  wire [4:0] ram_class_meta_field_type_14_field_type_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16]
  wire [2:0] ram_class_meta_field_type_14_field_type_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16]
  wire [4:0] ram_class_meta_field_type_14_field_type_MPORT_data; // @[Decoupled.scala 218:16]
  wire [2:0] ram_class_meta_field_type_14_field_type_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_class_meta_field_type_14_field_type_MPORT_mask; // @[Decoupled.scala 218:16]
  wire  ram_class_meta_field_type_14_field_type_MPORT_en; // @[Decoupled.scala 218:16]
  reg [15:0] ram_class_meta_field_type_14_sub_class_id [0:7]; // @[Decoupled.scala 218:16]
  wire [15:0] ram_class_meta_field_type_14_sub_class_id_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16]
  wire [2:0] ram_class_meta_field_type_14_sub_class_id_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16]
  wire [15:0] ram_class_meta_field_type_14_sub_class_id_MPORT_data; // @[Decoupled.scala 218:16]
  wire [2:0] ram_class_meta_field_type_14_sub_class_id_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_class_meta_field_type_14_sub_class_id_MPORT_mask; // @[Decoupled.scala 218:16]
  wire  ram_class_meta_field_type_14_sub_class_id_MPORT_en; // @[Decoupled.scala 218:16]
  reg  ram_class_meta_field_type_15_is_repeated [0:7]; // @[Decoupled.scala 218:16]
  wire  ram_class_meta_field_type_15_is_repeated_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16]
  wire [2:0] ram_class_meta_field_type_15_is_repeated_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_class_meta_field_type_15_is_repeated_MPORT_data; // @[Decoupled.scala 218:16]
  wire [2:0] ram_class_meta_field_type_15_is_repeated_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_class_meta_field_type_15_is_repeated_MPORT_mask; // @[Decoupled.scala 218:16]
  wire  ram_class_meta_field_type_15_is_repeated_MPORT_en; // @[Decoupled.scala 218:16]
  reg [4:0] ram_class_meta_field_type_15_field_type [0:7]; // @[Decoupled.scala 218:16]
  wire [4:0] ram_class_meta_field_type_15_field_type_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16]
  wire [2:0] ram_class_meta_field_type_15_field_type_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16]
  wire [4:0] ram_class_meta_field_type_15_field_type_MPORT_data; // @[Decoupled.scala 218:16]
  wire [2:0] ram_class_meta_field_type_15_field_type_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_class_meta_field_type_15_field_type_MPORT_mask; // @[Decoupled.scala 218:16]
  wire  ram_class_meta_field_type_15_field_type_MPORT_en; // @[Decoupled.scala 218:16]
  reg [15:0] ram_class_meta_field_type_15_sub_class_id [0:7]; // @[Decoupled.scala 218:16]
  wire [15:0] ram_class_meta_field_type_15_sub_class_id_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16]
  wire [2:0] ram_class_meta_field_type_15_sub_class_id_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16]
  wire [15:0] ram_class_meta_field_type_15_sub_class_id_MPORT_data; // @[Decoupled.scala 218:16]
  wire [2:0] ram_class_meta_field_type_15_sub_class_id_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_class_meta_field_type_15_sub_class_id_MPORT_mask; // @[Decoupled.scala 218:16]
  wire  ram_class_meta_field_type_15_sub_class_id_MPORT_en; // @[Decoupled.scala 218:16]
  reg  ram_class_meta_field_type_16_is_repeated [0:7]; // @[Decoupled.scala 218:16]
  wire  ram_class_meta_field_type_16_is_repeated_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16]
  wire [2:0] ram_class_meta_field_type_16_is_repeated_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_class_meta_field_type_16_is_repeated_MPORT_data; // @[Decoupled.scala 218:16]
  wire [2:0] ram_class_meta_field_type_16_is_repeated_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_class_meta_field_type_16_is_repeated_MPORT_mask; // @[Decoupled.scala 218:16]
  wire  ram_class_meta_field_type_16_is_repeated_MPORT_en; // @[Decoupled.scala 218:16]
  reg [4:0] ram_class_meta_field_type_16_field_type [0:7]; // @[Decoupled.scala 218:16]
  wire [4:0] ram_class_meta_field_type_16_field_type_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16]
  wire [2:0] ram_class_meta_field_type_16_field_type_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16]
  wire [4:0] ram_class_meta_field_type_16_field_type_MPORT_data; // @[Decoupled.scala 218:16]
  wire [2:0] ram_class_meta_field_type_16_field_type_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_class_meta_field_type_16_field_type_MPORT_mask; // @[Decoupled.scala 218:16]
  wire  ram_class_meta_field_type_16_field_type_MPORT_en; // @[Decoupled.scala 218:16]
  reg [15:0] ram_class_meta_field_type_16_sub_class_id [0:7]; // @[Decoupled.scala 218:16]
  wire [15:0] ram_class_meta_field_type_16_sub_class_id_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16]
  wire [2:0] ram_class_meta_field_type_16_sub_class_id_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16]
  wire [15:0] ram_class_meta_field_type_16_sub_class_id_MPORT_data; // @[Decoupled.scala 218:16]
  wire [2:0] ram_class_meta_field_type_16_sub_class_id_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_class_meta_field_type_16_sub_class_id_MPORT_mask; // @[Decoupled.scala 218:16]
  wire  ram_class_meta_field_type_16_sub_class_id_MPORT_en; // @[Decoupled.scala 218:16]
  reg  ram_class_meta_field_type_17_is_repeated [0:7]; // @[Decoupled.scala 218:16]
  wire  ram_class_meta_field_type_17_is_repeated_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16]
  wire [2:0] ram_class_meta_field_type_17_is_repeated_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_class_meta_field_type_17_is_repeated_MPORT_data; // @[Decoupled.scala 218:16]
  wire [2:0] ram_class_meta_field_type_17_is_repeated_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_class_meta_field_type_17_is_repeated_MPORT_mask; // @[Decoupled.scala 218:16]
  wire  ram_class_meta_field_type_17_is_repeated_MPORT_en; // @[Decoupled.scala 218:16]
  reg [4:0] ram_class_meta_field_type_17_field_type [0:7]; // @[Decoupled.scala 218:16]
  wire [4:0] ram_class_meta_field_type_17_field_type_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16]
  wire [2:0] ram_class_meta_field_type_17_field_type_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16]
  wire [4:0] ram_class_meta_field_type_17_field_type_MPORT_data; // @[Decoupled.scala 218:16]
  wire [2:0] ram_class_meta_field_type_17_field_type_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_class_meta_field_type_17_field_type_MPORT_mask; // @[Decoupled.scala 218:16]
  wire  ram_class_meta_field_type_17_field_type_MPORT_en; // @[Decoupled.scala 218:16]
  reg [15:0] ram_class_meta_field_type_17_sub_class_id [0:7]; // @[Decoupled.scala 218:16]
  wire [15:0] ram_class_meta_field_type_17_sub_class_id_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16]
  wire [2:0] ram_class_meta_field_type_17_sub_class_id_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16]
  wire [15:0] ram_class_meta_field_type_17_sub_class_id_MPORT_data; // @[Decoupled.scala 218:16]
  wire [2:0] ram_class_meta_field_type_17_sub_class_id_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_class_meta_field_type_17_sub_class_id_MPORT_mask; // @[Decoupled.scala 218:16]
  wire  ram_class_meta_field_type_17_sub_class_id_MPORT_en; // @[Decoupled.scala 218:16]
  reg  ram_class_meta_field_type_18_is_repeated [0:7]; // @[Decoupled.scala 218:16]
  wire  ram_class_meta_field_type_18_is_repeated_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16]
  wire [2:0] ram_class_meta_field_type_18_is_repeated_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_class_meta_field_type_18_is_repeated_MPORT_data; // @[Decoupled.scala 218:16]
  wire [2:0] ram_class_meta_field_type_18_is_repeated_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_class_meta_field_type_18_is_repeated_MPORT_mask; // @[Decoupled.scala 218:16]
  wire  ram_class_meta_field_type_18_is_repeated_MPORT_en; // @[Decoupled.scala 218:16]
  reg [4:0] ram_class_meta_field_type_18_field_type [0:7]; // @[Decoupled.scala 218:16]
  wire [4:0] ram_class_meta_field_type_18_field_type_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16]
  wire [2:0] ram_class_meta_field_type_18_field_type_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16]
  wire [4:0] ram_class_meta_field_type_18_field_type_MPORT_data; // @[Decoupled.scala 218:16]
  wire [2:0] ram_class_meta_field_type_18_field_type_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_class_meta_field_type_18_field_type_MPORT_mask; // @[Decoupled.scala 218:16]
  wire  ram_class_meta_field_type_18_field_type_MPORT_en; // @[Decoupled.scala 218:16]
  reg [15:0] ram_class_meta_field_type_18_sub_class_id [0:7]; // @[Decoupled.scala 218:16]
  wire [15:0] ram_class_meta_field_type_18_sub_class_id_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16]
  wire [2:0] ram_class_meta_field_type_18_sub_class_id_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16]
  wire [15:0] ram_class_meta_field_type_18_sub_class_id_MPORT_data; // @[Decoupled.scala 218:16]
  wire [2:0] ram_class_meta_field_type_18_sub_class_id_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_class_meta_field_type_18_sub_class_id_MPORT_mask; // @[Decoupled.scala 218:16]
  wire  ram_class_meta_field_type_18_sub_class_id_MPORT_en; // @[Decoupled.scala 218:16]
  reg  ram_class_meta_field_type_19_is_repeated [0:7]; // @[Decoupled.scala 218:16]
  wire  ram_class_meta_field_type_19_is_repeated_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16]
  wire [2:0] ram_class_meta_field_type_19_is_repeated_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_class_meta_field_type_19_is_repeated_MPORT_data; // @[Decoupled.scala 218:16]
  wire [2:0] ram_class_meta_field_type_19_is_repeated_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_class_meta_field_type_19_is_repeated_MPORT_mask; // @[Decoupled.scala 218:16]
  wire  ram_class_meta_field_type_19_is_repeated_MPORT_en; // @[Decoupled.scala 218:16]
  reg [4:0] ram_class_meta_field_type_19_field_type [0:7]; // @[Decoupled.scala 218:16]
  wire [4:0] ram_class_meta_field_type_19_field_type_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16]
  wire [2:0] ram_class_meta_field_type_19_field_type_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16]
  wire [4:0] ram_class_meta_field_type_19_field_type_MPORT_data; // @[Decoupled.scala 218:16]
  wire [2:0] ram_class_meta_field_type_19_field_type_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_class_meta_field_type_19_field_type_MPORT_mask; // @[Decoupled.scala 218:16]
  wire  ram_class_meta_field_type_19_field_type_MPORT_en; // @[Decoupled.scala 218:16]
  reg [15:0] ram_class_meta_field_type_19_sub_class_id [0:7]; // @[Decoupled.scala 218:16]
  wire [15:0] ram_class_meta_field_type_19_sub_class_id_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16]
  wire [2:0] ram_class_meta_field_type_19_sub_class_id_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16]
  wire [15:0] ram_class_meta_field_type_19_sub_class_id_MPORT_data; // @[Decoupled.scala 218:16]
  wire [2:0] ram_class_meta_field_type_19_sub_class_id_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_class_meta_field_type_19_sub_class_id_MPORT_mask; // @[Decoupled.scala 218:16]
  wire  ram_class_meta_field_type_19_sub_class_id_MPORT_en; // @[Decoupled.scala 218:16]
  reg  ram_class_meta_field_type_20_is_repeated [0:7]; // @[Decoupled.scala 218:16]
  wire  ram_class_meta_field_type_20_is_repeated_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16]
  wire [2:0] ram_class_meta_field_type_20_is_repeated_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_class_meta_field_type_20_is_repeated_MPORT_data; // @[Decoupled.scala 218:16]
  wire [2:0] ram_class_meta_field_type_20_is_repeated_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_class_meta_field_type_20_is_repeated_MPORT_mask; // @[Decoupled.scala 218:16]
  wire  ram_class_meta_field_type_20_is_repeated_MPORT_en; // @[Decoupled.scala 218:16]
  reg [4:0] ram_class_meta_field_type_20_field_type [0:7]; // @[Decoupled.scala 218:16]
  wire [4:0] ram_class_meta_field_type_20_field_type_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16]
  wire [2:0] ram_class_meta_field_type_20_field_type_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16]
  wire [4:0] ram_class_meta_field_type_20_field_type_MPORT_data; // @[Decoupled.scala 218:16]
  wire [2:0] ram_class_meta_field_type_20_field_type_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_class_meta_field_type_20_field_type_MPORT_mask; // @[Decoupled.scala 218:16]
  wire  ram_class_meta_field_type_20_field_type_MPORT_en; // @[Decoupled.scala 218:16]
  reg [15:0] ram_class_meta_field_type_20_sub_class_id [0:7]; // @[Decoupled.scala 218:16]
  wire [15:0] ram_class_meta_field_type_20_sub_class_id_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16]
  wire [2:0] ram_class_meta_field_type_20_sub_class_id_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16]
  wire [15:0] ram_class_meta_field_type_20_sub_class_id_MPORT_data; // @[Decoupled.scala 218:16]
  wire [2:0] ram_class_meta_field_type_20_sub_class_id_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_class_meta_field_type_20_sub_class_id_MPORT_mask; // @[Decoupled.scala 218:16]
  wire  ram_class_meta_field_type_20_sub_class_id_MPORT_en; // @[Decoupled.scala 218:16]
  reg  ram_class_meta_field_type_21_is_repeated [0:7]; // @[Decoupled.scala 218:16]
  wire  ram_class_meta_field_type_21_is_repeated_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16]
  wire [2:0] ram_class_meta_field_type_21_is_repeated_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_class_meta_field_type_21_is_repeated_MPORT_data; // @[Decoupled.scala 218:16]
  wire [2:0] ram_class_meta_field_type_21_is_repeated_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_class_meta_field_type_21_is_repeated_MPORT_mask; // @[Decoupled.scala 218:16]
  wire  ram_class_meta_field_type_21_is_repeated_MPORT_en; // @[Decoupled.scala 218:16]
  reg [4:0] ram_class_meta_field_type_21_field_type [0:7]; // @[Decoupled.scala 218:16]
  wire [4:0] ram_class_meta_field_type_21_field_type_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16]
  wire [2:0] ram_class_meta_field_type_21_field_type_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16]
  wire [4:0] ram_class_meta_field_type_21_field_type_MPORT_data; // @[Decoupled.scala 218:16]
  wire [2:0] ram_class_meta_field_type_21_field_type_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_class_meta_field_type_21_field_type_MPORT_mask; // @[Decoupled.scala 218:16]
  wire  ram_class_meta_field_type_21_field_type_MPORT_en; // @[Decoupled.scala 218:16]
  reg [15:0] ram_class_meta_field_type_21_sub_class_id [0:7]; // @[Decoupled.scala 218:16]
  wire [15:0] ram_class_meta_field_type_21_sub_class_id_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16]
  wire [2:0] ram_class_meta_field_type_21_sub_class_id_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16]
  wire [15:0] ram_class_meta_field_type_21_sub_class_id_MPORT_data; // @[Decoupled.scala 218:16]
  wire [2:0] ram_class_meta_field_type_21_sub_class_id_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_class_meta_field_type_21_sub_class_id_MPORT_mask; // @[Decoupled.scala 218:16]
  wire  ram_class_meta_field_type_21_sub_class_id_MPORT_en; // @[Decoupled.scala 218:16]
  reg  ram_class_meta_field_type_22_is_repeated [0:7]; // @[Decoupled.scala 218:16]
  wire  ram_class_meta_field_type_22_is_repeated_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16]
  wire [2:0] ram_class_meta_field_type_22_is_repeated_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_class_meta_field_type_22_is_repeated_MPORT_data; // @[Decoupled.scala 218:16]
  wire [2:0] ram_class_meta_field_type_22_is_repeated_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_class_meta_field_type_22_is_repeated_MPORT_mask; // @[Decoupled.scala 218:16]
  wire  ram_class_meta_field_type_22_is_repeated_MPORT_en; // @[Decoupled.scala 218:16]
  reg [4:0] ram_class_meta_field_type_22_field_type [0:7]; // @[Decoupled.scala 218:16]
  wire [4:0] ram_class_meta_field_type_22_field_type_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16]
  wire [2:0] ram_class_meta_field_type_22_field_type_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16]
  wire [4:0] ram_class_meta_field_type_22_field_type_MPORT_data; // @[Decoupled.scala 218:16]
  wire [2:0] ram_class_meta_field_type_22_field_type_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_class_meta_field_type_22_field_type_MPORT_mask; // @[Decoupled.scala 218:16]
  wire  ram_class_meta_field_type_22_field_type_MPORT_en; // @[Decoupled.scala 218:16]
  reg [15:0] ram_class_meta_field_type_22_sub_class_id [0:7]; // @[Decoupled.scala 218:16]
  wire [15:0] ram_class_meta_field_type_22_sub_class_id_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16]
  wire [2:0] ram_class_meta_field_type_22_sub_class_id_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16]
  wire [15:0] ram_class_meta_field_type_22_sub_class_id_MPORT_data; // @[Decoupled.scala 218:16]
  wire [2:0] ram_class_meta_field_type_22_sub_class_id_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_class_meta_field_type_22_sub_class_id_MPORT_mask; // @[Decoupled.scala 218:16]
  wire  ram_class_meta_field_type_22_sub_class_id_MPORT_en; // @[Decoupled.scala 218:16]
  reg  ram_class_meta_field_type_23_is_repeated [0:7]; // @[Decoupled.scala 218:16]
  wire  ram_class_meta_field_type_23_is_repeated_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16]
  wire [2:0] ram_class_meta_field_type_23_is_repeated_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_class_meta_field_type_23_is_repeated_MPORT_data; // @[Decoupled.scala 218:16]
  wire [2:0] ram_class_meta_field_type_23_is_repeated_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_class_meta_field_type_23_is_repeated_MPORT_mask; // @[Decoupled.scala 218:16]
  wire  ram_class_meta_field_type_23_is_repeated_MPORT_en; // @[Decoupled.scala 218:16]
  reg [4:0] ram_class_meta_field_type_23_field_type [0:7]; // @[Decoupled.scala 218:16]
  wire [4:0] ram_class_meta_field_type_23_field_type_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16]
  wire [2:0] ram_class_meta_field_type_23_field_type_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16]
  wire [4:0] ram_class_meta_field_type_23_field_type_MPORT_data; // @[Decoupled.scala 218:16]
  wire [2:0] ram_class_meta_field_type_23_field_type_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_class_meta_field_type_23_field_type_MPORT_mask; // @[Decoupled.scala 218:16]
  wire  ram_class_meta_field_type_23_field_type_MPORT_en; // @[Decoupled.scala 218:16]
  reg [15:0] ram_class_meta_field_type_23_sub_class_id [0:7]; // @[Decoupled.scala 218:16]
  wire [15:0] ram_class_meta_field_type_23_sub_class_id_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16]
  wire [2:0] ram_class_meta_field_type_23_sub_class_id_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16]
  wire [15:0] ram_class_meta_field_type_23_sub_class_id_MPORT_data; // @[Decoupled.scala 218:16]
  wire [2:0] ram_class_meta_field_type_23_sub_class_id_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_class_meta_field_type_23_sub_class_id_MPORT_mask; // @[Decoupled.scala 218:16]
  wire  ram_class_meta_field_type_23_sub_class_id_MPORT_en; // @[Decoupled.scala 218:16]
  reg  ram_class_meta_field_type_24_is_repeated [0:7]; // @[Decoupled.scala 218:16]
  wire  ram_class_meta_field_type_24_is_repeated_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16]
  wire [2:0] ram_class_meta_field_type_24_is_repeated_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_class_meta_field_type_24_is_repeated_MPORT_data; // @[Decoupled.scala 218:16]
  wire [2:0] ram_class_meta_field_type_24_is_repeated_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_class_meta_field_type_24_is_repeated_MPORT_mask; // @[Decoupled.scala 218:16]
  wire  ram_class_meta_field_type_24_is_repeated_MPORT_en; // @[Decoupled.scala 218:16]
  reg [4:0] ram_class_meta_field_type_24_field_type [0:7]; // @[Decoupled.scala 218:16]
  wire [4:0] ram_class_meta_field_type_24_field_type_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16]
  wire [2:0] ram_class_meta_field_type_24_field_type_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16]
  wire [4:0] ram_class_meta_field_type_24_field_type_MPORT_data; // @[Decoupled.scala 218:16]
  wire [2:0] ram_class_meta_field_type_24_field_type_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_class_meta_field_type_24_field_type_MPORT_mask; // @[Decoupled.scala 218:16]
  wire  ram_class_meta_field_type_24_field_type_MPORT_en; // @[Decoupled.scala 218:16]
  reg [15:0] ram_class_meta_field_type_24_sub_class_id [0:7]; // @[Decoupled.scala 218:16]
  wire [15:0] ram_class_meta_field_type_24_sub_class_id_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16]
  wire [2:0] ram_class_meta_field_type_24_sub_class_id_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16]
  wire [15:0] ram_class_meta_field_type_24_sub_class_id_MPORT_data; // @[Decoupled.scala 218:16]
  wire [2:0] ram_class_meta_field_type_24_sub_class_id_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_class_meta_field_type_24_sub_class_id_MPORT_mask; // @[Decoupled.scala 218:16]
  wire  ram_class_meta_field_type_24_sub_class_id_MPORT_en; // @[Decoupled.scala 218:16]
  reg  ram_class_meta_field_type_25_is_repeated [0:7]; // @[Decoupled.scala 218:16]
  wire  ram_class_meta_field_type_25_is_repeated_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16]
  wire [2:0] ram_class_meta_field_type_25_is_repeated_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_class_meta_field_type_25_is_repeated_MPORT_data; // @[Decoupled.scala 218:16]
  wire [2:0] ram_class_meta_field_type_25_is_repeated_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_class_meta_field_type_25_is_repeated_MPORT_mask; // @[Decoupled.scala 218:16]
  wire  ram_class_meta_field_type_25_is_repeated_MPORT_en; // @[Decoupled.scala 218:16]
  reg [4:0] ram_class_meta_field_type_25_field_type [0:7]; // @[Decoupled.scala 218:16]
  wire [4:0] ram_class_meta_field_type_25_field_type_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16]
  wire [2:0] ram_class_meta_field_type_25_field_type_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16]
  wire [4:0] ram_class_meta_field_type_25_field_type_MPORT_data; // @[Decoupled.scala 218:16]
  wire [2:0] ram_class_meta_field_type_25_field_type_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_class_meta_field_type_25_field_type_MPORT_mask; // @[Decoupled.scala 218:16]
  wire  ram_class_meta_field_type_25_field_type_MPORT_en; // @[Decoupled.scala 218:16]
  reg [15:0] ram_class_meta_field_type_25_sub_class_id [0:7]; // @[Decoupled.scala 218:16]
  wire [15:0] ram_class_meta_field_type_25_sub_class_id_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16]
  wire [2:0] ram_class_meta_field_type_25_sub_class_id_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16]
  wire [15:0] ram_class_meta_field_type_25_sub_class_id_MPORT_data; // @[Decoupled.scala 218:16]
  wire [2:0] ram_class_meta_field_type_25_sub_class_id_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_class_meta_field_type_25_sub_class_id_MPORT_mask; // @[Decoupled.scala 218:16]
  wire  ram_class_meta_field_type_25_sub_class_id_MPORT_en; // @[Decoupled.scala 218:16]
  reg  ram_class_meta_field_type_26_is_repeated [0:7]; // @[Decoupled.scala 218:16]
  wire  ram_class_meta_field_type_26_is_repeated_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16]
  wire [2:0] ram_class_meta_field_type_26_is_repeated_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_class_meta_field_type_26_is_repeated_MPORT_data; // @[Decoupled.scala 218:16]
  wire [2:0] ram_class_meta_field_type_26_is_repeated_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_class_meta_field_type_26_is_repeated_MPORT_mask; // @[Decoupled.scala 218:16]
  wire  ram_class_meta_field_type_26_is_repeated_MPORT_en; // @[Decoupled.scala 218:16]
  reg [4:0] ram_class_meta_field_type_26_field_type [0:7]; // @[Decoupled.scala 218:16]
  wire [4:0] ram_class_meta_field_type_26_field_type_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16]
  wire [2:0] ram_class_meta_field_type_26_field_type_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16]
  wire [4:0] ram_class_meta_field_type_26_field_type_MPORT_data; // @[Decoupled.scala 218:16]
  wire [2:0] ram_class_meta_field_type_26_field_type_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_class_meta_field_type_26_field_type_MPORT_mask; // @[Decoupled.scala 218:16]
  wire  ram_class_meta_field_type_26_field_type_MPORT_en; // @[Decoupled.scala 218:16]
  reg [15:0] ram_class_meta_field_type_26_sub_class_id [0:7]; // @[Decoupled.scala 218:16]
  wire [15:0] ram_class_meta_field_type_26_sub_class_id_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16]
  wire [2:0] ram_class_meta_field_type_26_sub_class_id_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16]
  wire [15:0] ram_class_meta_field_type_26_sub_class_id_MPORT_data; // @[Decoupled.scala 218:16]
  wire [2:0] ram_class_meta_field_type_26_sub_class_id_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_class_meta_field_type_26_sub_class_id_MPORT_mask; // @[Decoupled.scala 218:16]
  wire  ram_class_meta_field_type_26_sub_class_id_MPORT_en; // @[Decoupled.scala 218:16]
  reg  ram_class_meta_field_type_27_is_repeated [0:7]; // @[Decoupled.scala 218:16]
  wire  ram_class_meta_field_type_27_is_repeated_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16]
  wire [2:0] ram_class_meta_field_type_27_is_repeated_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_class_meta_field_type_27_is_repeated_MPORT_data; // @[Decoupled.scala 218:16]
  wire [2:0] ram_class_meta_field_type_27_is_repeated_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_class_meta_field_type_27_is_repeated_MPORT_mask; // @[Decoupled.scala 218:16]
  wire  ram_class_meta_field_type_27_is_repeated_MPORT_en; // @[Decoupled.scala 218:16]
  reg [4:0] ram_class_meta_field_type_27_field_type [0:7]; // @[Decoupled.scala 218:16]
  wire [4:0] ram_class_meta_field_type_27_field_type_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16]
  wire [2:0] ram_class_meta_field_type_27_field_type_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16]
  wire [4:0] ram_class_meta_field_type_27_field_type_MPORT_data; // @[Decoupled.scala 218:16]
  wire [2:0] ram_class_meta_field_type_27_field_type_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_class_meta_field_type_27_field_type_MPORT_mask; // @[Decoupled.scala 218:16]
  wire  ram_class_meta_field_type_27_field_type_MPORT_en; // @[Decoupled.scala 218:16]
  reg [15:0] ram_class_meta_field_type_27_sub_class_id [0:7]; // @[Decoupled.scala 218:16]
  wire [15:0] ram_class_meta_field_type_27_sub_class_id_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16]
  wire [2:0] ram_class_meta_field_type_27_sub_class_id_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16]
  wire [15:0] ram_class_meta_field_type_27_sub_class_id_MPORT_data; // @[Decoupled.scala 218:16]
  wire [2:0] ram_class_meta_field_type_27_sub_class_id_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_class_meta_field_type_27_sub_class_id_MPORT_mask; // @[Decoupled.scala 218:16]
  wire  ram_class_meta_field_type_27_sub_class_id_MPORT_en; // @[Decoupled.scala 218:16]
  reg  ram_class_meta_field_type_28_is_repeated [0:7]; // @[Decoupled.scala 218:16]
  wire  ram_class_meta_field_type_28_is_repeated_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16]
  wire [2:0] ram_class_meta_field_type_28_is_repeated_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_class_meta_field_type_28_is_repeated_MPORT_data; // @[Decoupled.scala 218:16]
  wire [2:0] ram_class_meta_field_type_28_is_repeated_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_class_meta_field_type_28_is_repeated_MPORT_mask; // @[Decoupled.scala 218:16]
  wire  ram_class_meta_field_type_28_is_repeated_MPORT_en; // @[Decoupled.scala 218:16]
  reg [4:0] ram_class_meta_field_type_28_field_type [0:7]; // @[Decoupled.scala 218:16]
  wire [4:0] ram_class_meta_field_type_28_field_type_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16]
  wire [2:0] ram_class_meta_field_type_28_field_type_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16]
  wire [4:0] ram_class_meta_field_type_28_field_type_MPORT_data; // @[Decoupled.scala 218:16]
  wire [2:0] ram_class_meta_field_type_28_field_type_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_class_meta_field_type_28_field_type_MPORT_mask; // @[Decoupled.scala 218:16]
  wire  ram_class_meta_field_type_28_field_type_MPORT_en; // @[Decoupled.scala 218:16]
  reg [15:0] ram_class_meta_field_type_28_sub_class_id [0:7]; // @[Decoupled.scala 218:16]
  wire [15:0] ram_class_meta_field_type_28_sub_class_id_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16]
  wire [2:0] ram_class_meta_field_type_28_sub_class_id_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16]
  wire [15:0] ram_class_meta_field_type_28_sub_class_id_MPORT_data; // @[Decoupled.scala 218:16]
  wire [2:0] ram_class_meta_field_type_28_sub_class_id_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_class_meta_field_type_28_sub_class_id_MPORT_mask; // @[Decoupled.scala 218:16]
  wire  ram_class_meta_field_type_28_sub_class_id_MPORT_en; // @[Decoupled.scala 218:16]
  reg  ram_class_meta_field_type_29_is_repeated [0:7]; // @[Decoupled.scala 218:16]
  wire  ram_class_meta_field_type_29_is_repeated_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16]
  wire [2:0] ram_class_meta_field_type_29_is_repeated_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_class_meta_field_type_29_is_repeated_MPORT_data; // @[Decoupled.scala 218:16]
  wire [2:0] ram_class_meta_field_type_29_is_repeated_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_class_meta_field_type_29_is_repeated_MPORT_mask; // @[Decoupled.scala 218:16]
  wire  ram_class_meta_field_type_29_is_repeated_MPORT_en; // @[Decoupled.scala 218:16]
  reg [4:0] ram_class_meta_field_type_29_field_type [0:7]; // @[Decoupled.scala 218:16]
  wire [4:0] ram_class_meta_field_type_29_field_type_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16]
  wire [2:0] ram_class_meta_field_type_29_field_type_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16]
  wire [4:0] ram_class_meta_field_type_29_field_type_MPORT_data; // @[Decoupled.scala 218:16]
  wire [2:0] ram_class_meta_field_type_29_field_type_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_class_meta_field_type_29_field_type_MPORT_mask; // @[Decoupled.scala 218:16]
  wire  ram_class_meta_field_type_29_field_type_MPORT_en; // @[Decoupled.scala 218:16]
  reg [15:0] ram_class_meta_field_type_29_sub_class_id [0:7]; // @[Decoupled.scala 218:16]
  wire [15:0] ram_class_meta_field_type_29_sub_class_id_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16]
  wire [2:0] ram_class_meta_field_type_29_sub_class_id_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16]
  wire [15:0] ram_class_meta_field_type_29_sub_class_id_MPORT_data; // @[Decoupled.scala 218:16]
  wire [2:0] ram_class_meta_field_type_29_sub_class_id_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_class_meta_field_type_29_sub_class_id_MPORT_mask; // @[Decoupled.scala 218:16]
  wire  ram_class_meta_field_type_29_sub_class_id_MPORT_en; // @[Decoupled.scala 218:16]
  reg  ram_class_meta_field_type_30_is_repeated [0:7]; // @[Decoupled.scala 218:16]
  wire  ram_class_meta_field_type_30_is_repeated_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16]
  wire [2:0] ram_class_meta_field_type_30_is_repeated_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_class_meta_field_type_30_is_repeated_MPORT_data; // @[Decoupled.scala 218:16]
  wire [2:0] ram_class_meta_field_type_30_is_repeated_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_class_meta_field_type_30_is_repeated_MPORT_mask; // @[Decoupled.scala 218:16]
  wire  ram_class_meta_field_type_30_is_repeated_MPORT_en; // @[Decoupled.scala 218:16]
  reg [4:0] ram_class_meta_field_type_30_field_type [0:7]; // @[Decoupled.scala 218:16]
  wire [4:0] ram_class_meta_field_type_30_field_type_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16]
  wire [2:0] ram_class_meta_field_type_30_field_type_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16]
  wire [4:0] ram_class_meta_field_type_30_field_type_MPORT_data; // @[Decoupled.scala 218:16]
  wire [2:0] ram_class_meta_field_type_30_field_type_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_class_meta_field_type_30_field_type_MPORT_mask; // @[Decoupled.scala 218:16]
  wire  ram_class_meta_field_type_30_field_type_MPORT_en; // @[Decoupled.scala 218:16]
  reg [15:0] ram_class_meta_field_type_30_sub_class_id [0:7]; // @[Decoupled.scala 218:16]
  wire [15:0] ram_class_meta_field_type_30_sub_class_id_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16]
  wire [2:0] ram_class_meta_field_type_30_sub_class_id_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16]
  wire [15:0] ram_class_meta_field_type_30_sub_class_id_MPORT_data; // @[Decoupled.scala 218:16]
  wire [2:0] ram_class_meta_field_type_30_sub_class_id_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_class_meta_field_type_30_sub_class_id_MPORT_mask; // @[Decoupled.scala 218:16]
  wire  ram_class_meta_field_type_30_sub_class_id_MPORT_en; // @[Decoupled.scala 218:16]
  reg  ram_class_meta_field_type_31_is_repeated [0:7]; // @[Decoupled.scala 218:16]
  wire  ram_class_meta_field_type_31_is_repeated_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16]
  wire [2:0] ram_class_meta_field_type_31_is_repeated_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_class_meta_field_type_31_is_repeated_MPORT_data; // @[Decoupled.scala 218:16]
  wire [2:0] ram_class_meta_field_type_31_is_repeated_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_class_meta_field_type_31_is_repeated_MPORT_mask; // @[Decoupled.scala 218:16]
  wire  ram_class_meta_field_type_31_is_repeated_MPORT_en; // @[Decoupled.scala 218:16]
  reg [4:0] ram_class_meta_field_type_31_field_type [0:7]; // @[Decoupled.scala 218:16]
  wire [4:0] ram_class_meta_field_type_31_field_type_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16]
  wire [2:0] ram_class_meta_field_type_31_field_type_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16]
  wire [4:0] ram_class_meta_field_type_31_field_type_MPORT_data; // @[Decoupled.scala 218:16]
  wire [2:0] ram_class_meta_field_type_31_field_type_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_class_meta_field_type_31_field_type_MPORT_mask; // @[Decoupled.scala 218:16]
  wire  ram_class_meta_field_type_31_field_type_MPORT_en; // @[Decoupled.scala 218:16]
  reg [15:0] ram_class_meta_field_type_31_sub_class_id [0:7]; // @[Decoupled.scala 218:16]
  wire [15:0] ram_class_meta_field_type_31_sub_class_id_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16]
  wire [2:0] ram_class_meta_field_type_31_sub_class_id_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16]
  wire [15:0] ram_class_meta_field_type_31_sub_class_id_MPORT_data; // @[Decoupled.scala 218:16]
  wire [2:0] ram_class_meta_field_type_31_sub_class_id_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_class_meta_field_type_31_sub_class_id_MPORT_mask; // @[Decoupled.scala 218:16]
  wire  ram_class_meta_field_type_31_sub_class_id_MPORT_en; // @[Decoupled.scala 218:16]
  reg  ram_class_meta_field_type_32_is_repeated [0:7]; // @[Decoupled.scala 218:16]
  wire  ram_class_meta_field_type_32_is_repeated_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16]
  wire [2:0] ram_class_meta_field_type_32_is_repeated_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_class_meta_field_type_32_is_repeated_MPORT_data; // @[Decoupled.scala 218:16]
  wire [2:0] ram_class_meta_field_type_32_is_repeated_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_class_meta_field_type_32_is_repeated_MPORT_mask; // @[Decoupled.scala 218:16]
  wire  ram_class_meta_field_type_32_is_repeated_MPORT_en; // @[Decoupled.scala 218:16]
  reg [4:0] ram_class_meta_field_type_32_field_type [0:7]; // @[Decoupled.scala 218:16]
  wire [4:0] ram_class_meta_field_type_32_field_type_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16]
  wire [2:0] ram_class_meta_field_type_32_field_type_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16]
  wire [4:0] ram_class_meta_field_type_32_field_type_MPORT_data; // @[Decoupled.scala 218:16]
  wire [2:0] ram_class_meta_field_type_32_field_type_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_class_meta_field_type_32_field_type_MPORT_mask; // @[Decoupled.scala 218:16]
  wire  ram_class_meta_field_type_32_field_type_MPORT_en; // @[Decoupled.scala 218:16]
  reg [15:0] ram_class_meta_field_type_32_sub_class_id [0:7]; // @[Decoupled.scala 218:16]
  wire [15:0] ram_class_meta_field_type_32_sub_class_id_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16]
  wire [2:0] ram_class_meta_field_type_32_sub_class_id_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16]
  wire [15:0] ram_class_meta_field_type_32_sub_class_id_MPORT_data; // @[Decoupled.scala 218:16]
  wire [2:0] ram_class_meta_field_type_32_sub_class_id_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_class_meta_field_type_32_sub_class_id_MPORT_mask; // @[Decoupled.scala 218:16]
  wire  ram_class_meta_field_type_32_sub_class_id_MPORT_en; // @[Decoupled.scala 218:16]
  reg [2:0] enq_ptr_value; // @[Counter.scala 60:40]
  reg [2:0] deq_ptr_value; // @[Counter.scala 60:40]
  reg  maybe_full; // @[Decoupled.scala 221:27]
  wire  ptr_match = enq_ptr_value == deq_ptr_value; // @[Decoupled.scala 223:33]
  wire  empty = ptr_match & ~maybe_full; // @[Decoupled.scala 224:25]
  wire  full = ptr_match & maybe_full; // @[Decoupled.scala 225:24]
  wire  do_enq = io_enq_ready & io_enq_valid; // @[Decoupled.scala 40:37]
  wire  do_deq = io_deq_ready & io_deq_valid; // @[Decoupled.scala 40:37]
  wire [2:0] _value_T_1 = enq_ptr_value + 3'h1; // @[Counter.scala 76:24]
  wire [2:0] _value_T_3 = deq_ptr_value + 3'h1; // @[Counter.scala 76:24]
  assign ram_class_meta_max_field_num_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_class_meta_max_field_num_io_deq_bits_MPORT_data =
    ram_class_meta_max_field_num[ram_class_meta_max_field_num_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  assign ram_class_meta_max_field_num_MPORT_data = io_enq_bits_class_meta_max_field_num;
  assign ram_class_meta_max_field_num_MPORT_addr = enq_ptr_value;
  assign ram_class_meta_max_field_num_MPORT_mask = 1'h1;
  assign ram_class_meta_max_field_num_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_class_meta_field_type_0_is_repeated_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_class_meta_field_type_0_is_repeated_io_deq_bits_MPORT_data =
    ram_class_meta_field_type_0_is_repeated[ram_class_meta_field_type_0_is_repeated_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  assign ram_class_meta_field_type_0_is_repeated_MPORT_data = io_enq_bits_class_meta_field_type_0_is_repeated;
  assign ram_class_meta_field_type_0_is_repeated_MPORT_addr = enq_ptr_value;
  assign ram_class_meta_field_type_0_is_repeated_MPORT_mask = 1'h1;
  assign ram_class_meta_field_type_0_is_repeated_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_class_meta_field_type_0_field_type_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_class_meta_field_type_0_field_type_io_deq_bits_MPORT_data =
    ram_class_meta_field_type_0_field_type[ram_class_meta_field_type_0_field_type_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  assign ram_class_meta_field_type_0_field_type_MPORT_data = io_enq_bits_class_meta_field_type_0_field_type;
  assign ram_class_meta_field_type_0_field_type_MPORT_addr = enq_ptr_value;
  assign ram_class_meta_field_type_0_field_type_MPORT_mask = 1'h1;
  assign ram_class_meta_field_type_0_field_type_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_class_meta_field_type_0_sub_class_id_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_class_meta_field_type_0_sub_class_id_io_deq_bits_MPORT_data =
    ram_class_meta_field_type_0_sub_class_id[ram_class_meta_field_type_0_sub_class_id_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  assign ram_class_meta_field_type_0_sub_class_id_MPORT_data = io_enq_bits_class_meta_field_type_0_sub_class_id;
  assign ram_class_meta_field_type_0_sub_class_id_MPORT_addr = enq_ptr_value;
  assign ram_class_meta_field_type_0_sub_class_id_MPORT_mask = 1'h1;
  assign ram_class_meta_field_type_0_sub_class_id_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_class_meta_field_type_1_is_repeated_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_class_meta_field_type_1_is_repeated_io_deq_bits_MPORT_data =
    ram_class_meta_field_type_1_is_repeated[ram_class_meta_field_type_1_is_repeated_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  assign ram_class_meta_field_type_1_is_repeated_MPORT_data = io_enq_bits_class_meta_field_type_1_is_repeated;
  assign ram_class_meta_field_type_1_is_repeated_MPORT_addr = enq_ptr_value;
  assign ram_class_meta_field_type_1_is_repeated_MPORT_mask = 1'h1;
  assign ram_class_meta_field_type_1_is_repeated_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_class_meta_field_type_1_field_type_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_class_meta_field_type_1_field_type_io_deq_bits_MPORT_data =
    ram_class_meta_field_type_1_field_type[ram_class_meta_field_type_1_field_type_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  assign ram_class_meta_field_type_1_field_type_MPORT_data = io_enq_bits_class_meta_field_type_1_field_type;
  assign ram_class_meta_field_type_1_field_type_MPORT_addr = enq_ptr_value;
  assign ram_class_meta_field_type_1_field_type_MPORT_mask = 1'h1;
  assign ram_class_meta_field_type_1_field_type_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_class_meta_field_type_1_sub_class_id_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_class_meta_field_type_1_sub_class_id_io_deq_bits_MPORT_data =
    ram_class_meta_field_type_1_sub_class_id[ram_class_meta_field_type_1_sub_class_id_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  assign ram_class_meta_field_type_1_sub_class_id_MPORT_data = io_enq_bits_class_meta_field_type_1_sub_class_id;
  assign ram_class_meta_field_type_1_sub_class_id_MPORT_addr = enq_ptr_value;
  assign ram_class_meta_field_type_1_sub_class_id_MPORT_mask = 1'h1;
  assign ram_class_meta_field_type_1_sub_class_id_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_class_meta_field_type_2_is_repeated_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_class_meta_field_type_2_is_repeated_io_deq_bits_MPORT_data =
    ram_class_meta_field_type_2_is_repeated[ram_class_meta_field_type_2_is_repeated_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  assign ram_class_meta_field_type_2_is_repeated_MPORT_data = io_enq_bits_class_meta_field_type_2_is_repeated;
  assign ram_class_meta_field_type_2_is_repeated_MPORT_addr = enq_ptr_value;
  assign ram_class_meta_field_type_2_is_repeated_MPORT_mask = 1'h1;
  assign ram_class_meta_field_type_2_is_repeated_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_class_meta_field_type_2_field_type_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_class_meta_field_type_2_field_type_io_deq_bits_MPORT_data =
    ram_class_meta_field_type_2_field_type[ram_class_meta_field_type_2_field_type_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  assign ram_class_meta_field_type_2_field_type_MPORT_data = io_enq_bits_class_meta_field_type_2_field_type;
  assign ram_class_meta_field_type_2_field_type_MPORT_addr = enq_ptr_value;
  assign ram_class_meta_field_type_2_field_type_MPORT_mask = 1'h1;
  assign ram_class_meta_field_type_2_field_type_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_class_meta_field_type_2_sub_class_id_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_class_meta_field_type_2_sub_class_id_io_deq_bits_MPORT_data =
    ram_class_meta_field_type_2_sub_class_id[ram_class_meta_field_type_2_sub_class_id_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  assign ram_class_meta_field_type_2_sub_class_id_MPORT_data = io_enq_bits_class_meta_field_type_2_sub_class_id;
  assign ram_class_meta_field_type_2_sub_class_id_MPORT_addr = enq_ptr_value;
  assign ram_class_meta_field_type_2_sub_class_id_MPORT_mask = 1'h1;
  assign ram_class_meta_field_type_2_sub_class_id_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_class_meta_field_type_3_is_repeated_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_class_meta_field_type_3_is_repeated_io_deq_bits_MPORT_data =
    ram_class_meta_field_type_3_is_repeated[ram_class_meta_field_type_3_is_repeated_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  assign ram_class_meta_field_type_3_is_repeated_MPORT_data = io_enq_bits_class_meta_field_type_3_is_repeated;
  assign ram_class_meta_field_type_3_is_repeated_MPORT_addr = enq_ptr_value;
  assign ram_class_meta_field_type_3_is_repeated_MPORT_mask = 1'h1;
  assign ram_class_meta_field_type_3_is_repeated_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_class_meta_field_type_3_field_type_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_class_meta_field_type_3_field_type_io_deq_bits_MPORT_data =
    ram_class_meta_field_type_3_field_type[ram_class_meta_field_type_3_field_type_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  assign ram_class_meta_field_type_3_field_type_MPORT_data = io_enq_bits_class_meta_field_type_3_field_type;
  assign ram_class_meta_field_type_3_field_type_MPORT_addr = enq_ptr_value;
  assign ram_class_meta_field_type_3_field_type_MPORT_mask = 1'h1;
  assign ram_class_meta_field_type_3_field_type_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_class_meta_field_type_3_sub_class_id_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_class_meta_field_type_3_sub_class_id_io_deq_bits_MPORT_data =
    ram_class_meta_field_type_3_sub_class_id[ram_class_meta_field_type_3_sub_class_id_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  assign ram_class_meta_field_type_3_sub_class_id_MPORT_data = io_enq_bits_class_meta_field_type_3_sub_class_id;
  assign ram_class_meta_field_type_3_sub_class_id_MPORT_addr = enq_ptr_value;
  assign ram_class_meta_field_type_3_sub_class_id_MPORT_mask = 1'h1;
  assign ram_class_meta_field_type_3_sub_class_id_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_class_meta_field_type_4_is_repeated_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_class_meta_field_type_4_is_repeated_io_deq_bits_MPORT_data =
    ram_class_meta_field_type_4_is_repeated[ram_class_meta_field_type_4_is_repeated_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  assign ram_class_meta_field_type_4_is_repeated_MPORT_data = io_enq_bits_class_meta_field_type_4_is_repeated;
  assign ram_class_meta_field_type_4_is_repeated_MPORT_addr = enq_ptr_value;
  assign ram_class_meta_field_type_4_is_repeated_MPORT_mask = 1'h1;
  assign ram_class_meta_field_type_4_is_repeated_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_class_meta_field_type_4_field_type_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_class_meta_field_type_4_field_type_io_deq_bits_MPORT_data =
    ram_class_meta_field_type_4_field_type[ram_class_meta_field_type_4_field_type_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  assign ram_class_meta_field_type_4_field_type_MPORT_data = io_enq_bits_class_meta_field_type_4_field_type;
  assign ram_class_meta_field_type_4_field_type_MPORT_addr = enq_ptr_value;
  assign ram_class_meta_field_type_4_field_type_MPORT_mask = 1'h1;
  assign ram_class_meta_field_type_4_field_type_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_class_meta_field_type_4_sub_class_id_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_class_meta_field_type_4_sub_class_id_io_deq_bits_MPORT_data =
    ram_class_meta_field_type_4_sub_class_id[ram_class_meta_field_type_4_sub_class_id_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  assign ram_class_meta_field_type_4_sub_class_id_MPORT_data = io_enq_bits_class_meta_field_type_4_sub_class_id;
  assign ram_class_meta_field_type_4_sub_class_id_MPORT_addr = enq_ptr_value;
  assign ram_class_meta_field_type_4_sub_class_id_MPORT_mask = 1'h1;
  assign ram_class_meta_field_type_4_sub_class_id_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_class_meta_field_type_5_is_repeated_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_class_meta_field_type_5_is_repeated_io_deq_bits_MPORT_data =
    ram_class_meta_field_type_5_is_repeated[ram_class_meta_field_type_5_is_repeated_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  assign ram_class_meta_field_type_5_is_repeated_MPORT_data = io_enq_bits_class_meta_field_type_5_is_repeated;
  assign ram_class_meta_field_type_5_is_repeated_MPORT_addr = enq_ptr_value;
  assign ram_class_meta_field_type_5_is_repeated_MPORT_mask = 1'h1;
  assign ram_class_meta_field_type_5_is_repeated_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_class_meta_field_type_5_field_type_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_class_meta_field_type_5_field_type_io_deq_bits_MPORT_data =
    ram_class_meta_field_type_5_field_type[ram_class_meta_field_type_5_field_type_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  assign ram_class_meta_field_type_5_field_type_MPORT_data = io_enq_bits_class_meta_field_type_5_field_type;
  assign ram_class_meta_field_type_5_field_type_MPORT_addr = enq_ptr_value;
  assign ram_class_meta_field_type_5_field_type_MPORT_mask = 1'h1;
  assign ram_class_meta_field_type_5_field_type_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_class_meta_field_type_5_sub_class_id_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_class_meta_field_type_5_sub_class_id_io_deq_bits_MPORT_data =
    ram_class_meta_field_type_5_sub_class_id[ram_class_meta_field_type_5_sub_class_id_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  assign ram_class_meta_field_type_5_sub_class_id_MPORT_data = io_enq_bits_class_meta_field_type_5_sub_class_id;
  assign ram_class_meta_field_type_5_sub_class_id_MPORT_addr = enq_ptr_value;
  assign ram_class_meta_field_type_5_sub_class_id_MPORT_mask = 1'h1;
  assign ram_class_meta_field_type_5_sub_class_id_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_class_meta_field_type_6_is_repeated_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_class_meta_field_type_6_is_repeated_io_deq_bits_MPORT_data =
    ram_class_meta_field_type_6_is_repeated[ram_class_meta_field_type_6_is_repeated_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  assign ram_class_meta_field_type_6_is_repeated_MPORT_data = io_enq_bits_class_meta_field_type_6_is_repeated;
  assign ram_class_meta_field_type_6_is_repeated_MPORT_addr = enq_ptr_value;
  assign ram_class_meta_field_type_6_is_repeated_MPORT_mask = 1'h1;
  assign ram_class_meta_field_type_6_is_repeated_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_class_meta_field_type_6_field_type_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_class_meta_field_type_6_field_type_io_deq_bits_MPORT_data =
    ram_class_meta_field_type_6_field_type[ram_class_meta_field_type_6_field_type_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  assign ram_class_meta_field_type_6_field_type_MPORT_data = io_enq_bits_class_meta_field_type_6_field_type;
  assign ram_class_meta_field_type_6_field_type_MPORT_addr = enq_ptr_value;
  assign ram_class_meta_field_type_6_field_type_MPORT_mask = 1'h1;
  assign ram_class_meta_field_type_6_field_type_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_class_meta_field_type_6_sub_class_id_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_class_meta_field_type_6_sub_class_id_io_deq_bits_MPORT_data =
    ram_class_meta_field_type_6_sub_class_id[ram_class_meta_field_type_6_sub_class_id_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  assign ram_class_meta_field_type_6_sub_class_id_MPORT_data = io_enq_bits_class_meta_field_type_6_sub_class_id;
  assign ram_class_meta_field_type_6_sub_class_id_MPORT_addr = enq_ptr_value;
  assign ram_class_meta_field_type_6_sub_class_id_MPORT_mask = 1'h1;
  assign ram_class_meta_field_type_6_sub_class_id_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_class_meta_field_type_7_is_repeated_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_class_meta_field_type_7_is_repeated_io_deq_bits_MPORT_data =
    ram_class_meta_field_type_7_is_repeated[ram_class_meta_field_type_7_is_repeated_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  assign ram_class_meta_field_type_7_is_repeated_MPORT_data = io_enq_bits_class_meta_field_type_7_is_repeated;
  assign ram_class_meta_field_type_7_is_repeated_MPORT_addr = enq_ptr_value;
  assign ram_class_meta_field_type_7_is_repeated_MPORT_mask = 1'h1;
  assign ram_class_meta_field_type_7_is_repeated_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_class_meta_field_type_7_field_type_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_class_meta_field_type_7_field_type_io_deq_bits_MPORT_data =
    ram_class_meta_field_type_7_field_type[ram_class_meta_field_type_7_field_type_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  assign ram_class_meta_field_type_7_field_type_MPORT_data = io_enq_bits_class_meta_field_type_7_field_type;
  assign ram_class_meta_field_type_7_field_type_MPORT_addr = enq_ptr_value;
  assign ram_class_meta_field_type_7_field_type_MPORT_mask = 1'h1;
  assign ram_class_meta_field_type_7_field_type_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_class_meta_field_type_7_sub_class_id_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_class_meta_field_type_7_sub_class_id_io_deq_bits_MPORT_data =
    ram_class_meta_field_type_7_sub_class_id[ram_class_meta_field_type_7_sub_class_id_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  assign ram_class_meta_field_type_7_sub_class_id_MPORT_data = io_enq_bits_class_meta_field_type_7_sub_class_id;
  assign ram_class_meta_field_type_7_sub_class_id_MPORT_addr = enq_ptr_value;
  assign ram_class_meta_field_type_7_sub_class_id_MPORT_mask = 1'h1;
  assign ram_class_meta_field_type_7_sub_class_id_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_class_meta_field_type_8_is_repeated_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_class_meta_field_type_8_is_repeated_io_deq_bits_MPORT_data =
    ram_class_meta_field_type_8_is_repeated[ram_class_meta_field_type_8_is_repeated_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  assign ram_class_meta_field_type_8_is_repeated_MPORT_data = io_enq_bits_class_meta_field_type_8_is_repeated;
  assign ram_class_meta_field_type_8_is_repeated_MPORT_addr = enq_ptr_value;
  assign ram_class_meta_field_type_8_is_repeated_MPORT_mask = 1'h1;
  assign ram_class_meta_field_type_8_is_repeated_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_class_meta_field_type_8_field_type_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_class_meta_field_type_8_field_type_io_deq_bits_MPORT_data =
    ram_class_meta_field_type_8_field_type[ram_class_meta_field_type_8_field_type_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  assign ram_class_meta_field_type_8_field_type_MPORT_data = io_enq_bits_class_meta_field_type_8_field_type;
  assign ram_class_meta_field_type_8_field_type_MPORT_addr = enq_ptr_value;
  assign ram_class_meta_field_type_8_field_type_MPORT_mask = 1'h1;
  assign ram_class_meta_field_type_8_field_type_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_class_meta_field_type_8_sub_class_id_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_class_meta_field_type_8_sub_class_id_io_deq_bits_MPORT_data =
    ram_class_meta_field_type_8_sub_class_id[ram_class_meta_field_type_8_sub_class_id_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  assign ram_class_meta_field_type_8_sub_class_id_MPORT_data = io_enq_bits_class_meta_field_type_8_sub_class_id;
  assign ram_class_meta_field_type_8_sub_class_id_MPORT_addr = enq_ptr_value;
  assign ram_class_meta_field_type_8_sub_class_id_MPORT_mask = 1'h1;
  assign ram_class_meta_field_type_8_sub_class_id_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_class_meta_field_type_9_is_repeated_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_class_meta_field_type_9_is_repeated_io_deq_bits_MPORT_data =
    ram_class_meta_field_type_9_is_repeated[ram_class_meta_field_type_9_is_repeated_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  assign ram_class_meta_field_type_9_is_repeated_MPORT_data = io_enq_bits_class_meta_field_type_9_is_repeated;
  assign ram_class_meta_field_type_9_is_repeated_MPORT_addr = enq_ptr_value;
  assign ram_class_meta_field_type_9_is_repeated_MPORT_mask = 1'h1;
  assign ram_class_meta_field_type_9_is_repeated_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_class_meta_field_type_9_field_type_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_class_meta_field_type_9_field_type_io_deq_bits_MPORT_data =
    ram_class_meta_field_type_9_field_type[ram_class_meta_field_type_9_field_type_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  assign ram_class_meta_field_type_9_field_type_MPORT_data = io_enq_bits_class_meta_field_type_9_field_type;
  assign ram_class_meta_field_type_9_field_type_MPORT_addr = enq_ptr_value;
  assign ram_class_meta_field_type_9_field_type_MPORT_mask = 1'h1;
  assign ram_class_meta_field_type_9_field_type_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_class_meta_field_type_9_sub_class_id_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_class_meta_field_type_9_sub_class_id_io_deq_bits_MPORT_data =
    ram_class_meta_field_type_9_sub_class_id[ram_class_meta_field_type_9_sub_class_id_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  assign ram_class_meta_field_type_9_sub_class_id_MPORT_data = io_enq_bits_class_meta_field_type_9_sub_class_id;
  assign ram_class_meta_field_type_9_sub_class_id_MPORT_addr = enq_ptr_value;
  assign ram_class_meta_field_type_9_sub_class_id_MPORT_mask = 1'h1;
  assign ram_class_meta_field_type_9_sub_class_id_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_class_meta_field_type_10_is_repeated_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_class_meta_field_type_10_is_repeated_io_deq_bits_MPORT_data =
    ram_class_meta_field_type_10_is_repeated[ram_class_meta_field_type_10_is_repeated_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  assign ram_class_meta_field_type_10_is_repeated_MPORT_data = io_enq_bits_class_meta_field_type_10_is_repeated;
  assign ram_class_meta_field_type_10_is_repeated_MPORT_addr = enq_ptr_value;
  assign ram_class_meta_field_type_10_is_repeated_MPORT_mask = 1'h1;
  assign ram_class_meta_field_type_10_is_repeated_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_class_meta_field_type_10_field_type_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_class_meta_field_type_10_field_type_io_deq_bits_MPORT_data =
    ram_class_meta_field_type_10_field_type[ram_class_meta_field_type_10_field_type_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  assign ram_class_meta_field_type_10_field_type_MPORT_data = io_enq_bits_class_meta_field_type_10_field_type;
  assign ram_class_meta_field_type_10_field_type_MPORT_addr = enq_ptr_value;
  assign ram_class_meta_field_type_10_field_type_MPORT_mask = 1'h1;
  assign ram_class_meta_field_type_10_field_type_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_class_meta_field_type_10_sub_class_id_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_class_meta_field_type_10_sub_class_id_io_deq_bits_MPORT_data =
    ram_class_meta_field_type_10_sub_class_id[ram_class_meta_field_type_10_sub_class_id_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  assign ram_class_meta_field_type_10_sub_class_id_MPORT_data = io_enq_bits_class_meta_field_type_10_sub_class_id;
  assign ram_class_meta_field_type_10_sub_class_id_MPORT_addr = enq_ptr_value;
  assign ram_class_meta_field_type_10_sub_class_id_MPORT_mask = 1'h1;
  assign ram_class_meta_field_type_10_sub_class_id_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_class_meta_field_type_11_is_repeated_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_class_meta_field_type_11_is_repeated_io_deq_bits_MPORT_data =
    ram_class_meta_field_type_11_is_repeated[ram_class_meta_field_type_11_is_repeated_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  assign ram_class_meta_field_type_11_is_repeated_MPORT_data = io_enq_bits_class_meta_field_type_11_is_repeated;
  assign ram_class_meta_field_type_11_is_repeated_MPORT_addr = enq_ptr_value;
  assign ram_class_meta_field_type_11_is_repeated_MPORT_mask = 1'h1;
  assign ram_class_meta_field_type_11_is_repeated_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_class_meta_field_type_11_field_type_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_class_meta_field_type_11_field_type_io_deq_bits_MPORT_data =
    ram_class_meta_field_type_11_field_type[ram_class_meta_field_type_11_field_type_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  assign ram_class_meta_field_type_11_field_type_MPORT_data = io_enq_bits_class_meta_field_type_11_field_type;
  assign ram_class_meta_field_type_11_field_type_MPORT_addr = enq_ptr_value;
  assign ram_class_meta_field_type_11_field_type_MPORT_mask = 1'h1;
  assign ram_class_meta_field_type_11_field_type_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_class_meta_field_type_11_sub_class_id_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_class_meta_field_type_11_sub_class_id_io_deq_bits_MPORT_data =
    ram_class_meta_field_type_11_sub_class_id[ram_class_meta_field_type_11_sub_class_id_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  assign ram_class_meta_field_type_11_sub_class_id_MPORT_data = io_enq_bits_class_meta_field_type_11_sub_class_id;
  assign ram_class_meta_field_type_11_sub_class_id_MPORT_addr = enq_ptr_value;
  assign ram_class_meta_field_type_11_sub_class_id_MPORT_mask = 1'h1;
  assign ram_class_meta_field_type_11_sub_class_id_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_class_meta_field_type_12_is_repeated_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_class_meta_field_type_12_is_repeated_io_deq_bits_MPORT_data =
    ram_class_meta_field_type_12_is_repeated[ram_class_meta_field_type_12_is_repeated_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  assign ram_class_meta_field_type_12_is_repeated_MPORT_data = io_enq_bits_class_meta_field_type_12_is_repeated;
  assign ram_class_meta_field_type_12_is_repeated_MPORT_addr = enq_ptr_value;
  assign ram_class_meta_field_type_12_is_repeated_MPORT_mask = 1'h1;
  assign ram_class_meta_field_type_12_is_repeated_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_class_meta_field_type_12_field_type_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_class_meta_field_type_12_field_type_io_deq_bits_MPORT_data =
    ram_class_meta_field_type_12_field_type[ram_class_meta_field_type_12_field_type_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  assign ram_class_meta_field_type_12_field_type_MPORT_data = io_enq_bits_class_meta_field_type_12_field_type;
  assign ram_class_meta_field_type_12_field_type_MPORT_addr = enq_ptr_value;
  assign ram_class_meta_field_type_12_field_type_MPORT_mask = 1'h1;
  assign ram_class_meta_field_type_12_field_type_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_class_meta_field_type_12_sub_class_id_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_class_meta_field_type_12_sub_class_id_io_deq_bits_MPORT_data =
    ram_class_meta_field_type_12_sub_class_id[ram_class_meta_field_type_12_sub_class_id_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  assign ram_class_meta_field_type_12_sub_class_id_MPORT_data = io_enq_bits_class_meta_field_type_12_sub_class_id;
  assign ram_class_meta_field_type_12_sub_class_id_MPORT_addr = enq_ptr_value;
  assign ram_class_meta_field_type_12_sub_class_id_MPORT_mask = 1'h1;
  assign ram_class_meta_field_type_12_sub_class_id_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_class_meta_field_type_13_is_repeated_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_class_meta_field_type_13_is_repeated_io_deq_bits_MPORT_data =
    ram_class_meta_field_type_13_is_repeated[ram_class_meta_field_type_13_is_repeated_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  assign ram_class_meta_field_type_13_is_repeated_MPORT_data = io_enq_bits_class_meta_field_type_13_is_repeated;
  assign ram_class_meta_field_type_13_is_repeated_MPORT_addr = enq_ptr_value;
  assign ram_class_meta_field_type_13_is_repeated_MPORT_mask = 1'h1;
  assign ram_class_meta_field_type_13_is_repeated_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_class_meta_field_type_13_field_type_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_class_meta_field_type_13_field_type_io_deq_bits_MPORT_data =
    ram_class_meta_field_type_13_field_type[ram_class_meta_field_type_13_field_type_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  assign ram_class_meta_field_type_13_field_type_MPORT_data = io_enq_bits_class_meta_field_type_13_field_type;
  assign ram_class_meta_field_type_13_field_type_MPORT_addr = enq_ptr_value;
  assign ram_class_meta_field_type_13_field_type_MPORT_mask = 1'h1;
  assign ram_class_meta_field_type_13_field_type_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_class_meta_field_type_13_sub_class_id_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_class_meta_field_type_13_sub_class_id_io_deq_bits_MPORT_data =
    ram_class_meta_field_type_13_sub_class_id[ram_class_meta_field_type_13_sub_class_id_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  assign ram_class_meta_field_type_13_sub_class_id_MPORT_data = io_enq_bits_class_meta_field_type_13_sub_class_id;
  assign ram_class_meta_field_type_13_sub_class_id_MPORT_addr = enq_ptr_value;
  assign ram_class_meta_field_type_13_sub_class_id_MPORT_mask = 1'h1;
  assign ram_class_meta_field_type_13_sub_class_id_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_class_meta_field_type_14_is_repeated_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_class_meta_field_type_14_is_repeated_io_deq_bits_MPORT_data =
    ram_class_meta_field_type_14_is_repeated[ram_class_meta_field_type_14_is_repeated_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  assign ram_class_meta_field_type_14_is_repeated_MPORT_data = io_enq_bits_class_meta_field_type_14_is_repeated;
  assign ram_class_meta_field_type_14_is_repeated_MPORT_addr = enq_ptr_value;
  assign ram_class_meta_field_type_14_is_repeated_MPORT_mask = 1'h1;
  assign ram_class_meta_field_type_14_is_repeated_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_class_meta_field_type_14_field_type_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_class_meta_field_type_14_field_type_io_deq_bits_MPORT_data =
    ram_class_meta_field_type_14_field_type[ram_class_meta_field_type_14_field_type_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  assign ram_class_meta_field_type_14_field_type_MPORT_data = io_enq_bits_class_meta_field_type_14_field_type;
  assign ram_class_meta_field_type_14_field_type_MPORT_addr = enq_ptr_value;
  assign ram_class_meta_field_type_14_field_type_MPORT_mask = 1'h1;
  assign ram_class_meta_field_type_14_field_type_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_class_meta_field_type_14_sub_class_id_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_class_meta_field_type_14_sub_class_id_io_deq_bits_MPORT_data =
    ram_class_meta_field_type_14_sub_class_id[ram_class_meta_field_type_14_sub_class_id_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  assign ram_class_meta_field_type_14_sub_class_id_MPORT_data = io_enq_bits_class_meta_field_type_14_sub_class_id;
  assign ram_class_meta_field_type_14_sub_class_id_MPORT_addr = enq_ptr_value;
  assign ram_class_meta_field_type_14_sub_class_id_MPORT_mask = 1'h1;
  assign ram_class_meta_field_type_14_sub_class_id_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_class_meta_field_type_15_is_repeated_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_class_meta_field_type_15_is_repeated_io_deq_bits_MPORT_data =
    ram_class_meta_field_type_15_is_repeated[ram_class_meta_field_type_15_is_repeated_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  assign ram_class_meta_field_type_15_is_repeated_MPORT_data = io_enq_bits_class_meta_field_type_15_is_repeated;
  assign ram_class_meta_field_type_15_is_repeated_MPORT_addr = enq_ptr_value;
  assign ram_class_meta_field_type_15_is_repeated_MPORT_mask = 1'h1;
  assign ram_class_meta_field_type_15_is_repeated_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_class_meta_field_type_15_field_type_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_class_meta_field_type_15_field_type_io_deq_bits_MPORT_data =
    ram_class_meta_field_type_15_field_type[ram_class_meta_field_type_15_field_type_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  assign ram_class_meta_field_type_15_field_type_MPORT_data = io_enq_bits_class_meta_field_type_15_field_type;
  assign ram_class_meta_field_type_15_field_type_MPORT_addr = enq_ptr_value;
  assign ram_class_meta_field_type_15_field_type_MPORT_mask = 1'h1;
  assign ram_class_meta_field_type_15_field_type_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_class_meta_field_type_15_sub_class_id_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_class_meta_field_type_15_sub_class_id_io_deq_bits_MPORT_data =
    ram_class_meta_field_type_15_sub_class_id[ram_class_meta_field_type_15_sub_class_id_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  assign ram_class_meta_field_type_15_sub_class_id_MPORT_data = io_enq_bits_class_meta_field_type_15_sub_class_id;
  assign ram_class_meta_field_type_15_sub_class_id_MPORT_addr = enq_ptr_value;
  assign ram_class_meta_field_type_15_sub_class_id_MPORT_mask = 1'h1;
  assign ram_class_meta_field_type_15_sub_class_id_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_class_meta_field_type_16_is_repeated_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_class_meta_field_type_16_is_repeated_io_deq_bits_MPORT_data =
    ram_class_meta_field_type_16_is_repeated[ram_class_meta_field_type_16_is_repeated_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  assign ram_class_meta_field_type_16_is_repeated_MPORT_data = io_enq_bits_class_meta_field_type_16_is_repeated;
  assign ram_class_meta_field_type_16_is_repeated_MPORT_addr = enq_ptr_value;
  assign ram_class_meta_field_type_16_is_repeated_MPORT_mask = 1'h1;
  assign ram_class_meta_field_type_16_is_repeated_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_class_meta_field_type_16_field_type_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_class_meta_field_type_16_field_type_io_deq_bits_MPORT_data =
    ram_class_meta_field_type_16_field_type[ram_class_meta_field_type_16_field_type_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  assign ram_class_meta_field_type_16_field_type_MPORT_data = io_enq_bits_class_meta_field_type_16_field_type;
  assign ram_class_meta_field_type_16_field_type_MPORT_addr = enq_ptr_value;
  assign ram_class_meta_field_type_16_field_type_MPORT_mask = 1'h1;
  assign ram_class_meta_field_type_16_field_type_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_class_meta_field_type_16_sub_class_id_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_class_meta_field_type_16_sub_class_id_io_deq_bits_MPORT_data =
    ram_class_meta_field_type_16_sub_class_id[ram_class_meta_field_type_16_sub_class_id_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  assign ram_class_meta_field_type_16_sub_class_id_MPORT_data = io_enq_bits_class_meta_field_type_16_sub_class_id;
  assign ram_class_meta_field_type_16_sub_class_id_MPORT_addr = enq_ptr_value;
  assign ram_class_meta_field_type_16_sub_class_id_MPORT_mask = 1'h1;
  assign ram_class_meta_field_type_16_sub_class_id_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_class_meta_field_type_17_is_repeated_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_class_meta_field_type_17_is_repeated_io_deq_bits_MPORT_data =
    ram_class_meta_field_type_17_is_repeated[ram_class_meta_field_type_17_is_repeated_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  assign ram_class_meta_field_type_17_is_repeated_MPORT_data = io_enq_bits_class_meta_field_type_17_is_repeated;
  assign ram_class_meta_field_type_17_is_repeated_MPORT_addr = enq_ptr_value;
  assign ram_class_meta_field_type_17_is_repeated_MPORT_mask = 1'h1;
  assign ram_class_meta_field_type_17_is_repeated_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_class_meta_field_type_17_field_type_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_class_meta_field_type_17_field_type_io_deq_bits_MPORT_data =
    ram_class_meta_field_type_17_field_type[ram_class_meta_field_type_17_field_type_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  assign ram_class_meta_field_type_17_field_type_MPORT_data = io_enq_bits_class_meta_field_type_17_field_type;
  assign ram_class_meta_field_type_17_field_type_MPORT_addr = enq_ptr_value;
  assign ram_class_meta_field_type_17_field_type_MPORT_mask = 1'h1;
  assign ram_class_meta_field_type_17_field_type_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_class_meta_field_type_17_sub_class_id_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_class_meta_field_type_17_sub_class_id_io_deq_bits_MPORT_data =
    ram_class_meta_field_type_17_sub_class_id[ram_class_meta_field_type_17_sub_class_id_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  assign ram_class_meta_field_type_17_sub_class_id_MPORT_data = io_enq_bits_class_meta_field_type_17_sub_class_id;
  assign ram_class_meta_field_type_17_sub_class_id_MPORT_addr = enq_ptr_value;
  assign ram_class_meta_field_type_17_sub_class_id_MPORT_mask = 1'h1;
  assign ram_class_meta_field_type_17_sub_class_id_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_class_meta_field_type_18_is_repeated_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_class_meta_field_type_18_is_repeated_io_deq_bits_MPORT_data =
    ram_class_meta_field_type_18_is_repeated[ram_class_meta_field_type_18_is_repeated_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  assign ram_class_meta_field_type_18_is_repeated_MPORT_data = io_enq_bits_class_meta_field_type_18_is_repeated;
  assign ram_class_meta_field_type_18_is_repeated_MPORT_addr = enq_ptr_value;
  assign ram_class_meta_field_type_18_is_repeated_MPORT_mask = 1'h1;
  assign ram_class_meta_field_type_18_is_repeated_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_class_meta_field_type_18_field_type_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_class_meta_field_type_18_field_type_io_deq_bits_MPORT_data =
    ram_class_meta_field_type_18_field_type[ram_class_meta_field_type_18_field_type_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  assign ram_class_meta_field_type_18_field_type_MPORT_data = io_enq_bits_class_meta_field_type_18_field_type;
  assign ram_class_meta_field_type_18_field_type_MPORT_addr = enq_ptr_value;
  assign ram_class_meta_field_type_18_field_type_MPORT_mask = 1'h1;
  assign ram_class_meta_field_type_18_field_type_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_class_meta_field_type_18_sub_class_id_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_class_meta_field_type_18_sub_class_id_io_deq_bits_MPORT_data =
    ram_class_meta_field_type_18_sub_class_id[ram_class_meta_field_type_18_sub_class_id_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  assign ram_class_meta_field_type_18_sub_class_id_MPORT_data = io_enq_bits_class_meta_field_type_18_sub_class_id;
  assign ram_class_meta_field_type_18_sub_class_id_MPORT_addr = enq_ptr_value;
  assign ram_class_meta_field_type_18_sub_class_id_MPORT_mask = 1'h1;
  assign ram_class_meta_field_type_18_sub_class_id_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_class_meta_field_type_19_is_repeated_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_class_meta_field_type_19_is_repeated_io_deq_bits_MPORT_data =
    ram_class_meta_field_type_19_is_repeated[ram_class_meta_field_type_19_is_repeated_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  assign ram_class_meta_field_type_19_is_repeated_MPORT_data = io_enq_bits_class_meta_field_type_19_is_repeated;
  assign ram_class_meta_field_type_19_is_repeated_MPORT_addr = enq_ptr_value;
  assign ram_class_meta_field_type_19_is_repeated_MPORT_mask = 1'h1;
  assign ram_class_meta_field_type_19_is_repeated_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_class_meta_field_type_19_field_type_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_class_meta_field_type_19_field_type_io_deq_bits_MPORT_data =
    ram_class_meta_field_type_19_field_type[ram_class_meta_field_type_19_field_type_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  assign ram_class_meta_field_type_19_field_type_MPORT_data = io_enq_bits_class_meta_field_type_19_field_type;
  assign ram_class_meta_field_type_19_field_type_MPORT_addr = enq_ptr_value;
  assign ram_class_meta_field_type_19_field_type_MPORT_mask = 1'h1;
  assign ram_class_meta_field_type_19_field_type_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_class_meta_field_type_19_sub_class_id_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_class_meta_field_type_19_sub_class_id_io_deq_bits_MPORT_data =
    ram_class_meta_field_type_19_sub_class_id[ram_class_meta_field_type_19_sub_class_id_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  assign ram_class_meta_field_type_19_sub_class_id_MPORT_data = io_enq_bits_class_meta_field_type_19_sub_class_id;
  assign ram_class_meta_field_type_19_sub_class_id_MPORT_addr = enq_ptr_value;
  assign ram_class_meta_field_type_19_sub_class_id_MPORT_mask = 1'h1;
  assign ram_class_meta_field_type_19_sub_class_id_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_class_meta_field_type_20_is_repeated_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_class_meta_field_type_20_is_repeated_io_deq_bits_MPORT_data =
    ram_class_meta_field_type_20_is_repeated[ram_class_meta_field_type_20_is_repeated_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  assign ram_class_meta_field_type_20_is_repeated_MPORT_data = io_enq_bits_class_meta_field_type_20_is_repeated;
  assign ram_class_meta_field_type_20_is_repeated_MPORT_addr = enq_ptr_value;
  assign ram_class_meta_field_type_20_is_repeated_MPORT_mask = 1'h1;
  assign ram_class_meta_field_type_20_is_repeated_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_class_meta_field_type_20_field_type_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_class_meta_field_type_20_field_type_io_deq_bits_MPORT_data =
    ram_class_meta_field_type_20_field_type[ram_class_meta_field_type_20_field_type_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  assign ram_class_meta_field_type_20_field_type_MPORT_data = io_enq_bits_class_meta_field_type_20_field_type;
  assign ram_class_meta_field_type_20_field_type_MPORT_addr = enq_ptr_value;
  assign ram_class_meta_field_type_20_field_type_MPORT_mask = 1'h1;
  assign ram_class_meta_field_type_20_field_type_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_class_meta_field_type_20_sub_class_id_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_class_meta_field_type_20_sub_class_id_io_deq_bits_MPORT_data =
    ram_class_meta_field_type_20_sub_class_id[ram_class_meta_field_type_20_sub_class_id_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  assign ram_class_meta_field_type_20_sub_class_id_MPORT_data = io_enq_bits_class_meta_field_type_20_sub_class_id;
  assign ram_class_meta_field_type_20_sub_class_id_MPORT_addr = enq_ptr_value;
  assign ram_class_meta_field_type_20_sub_class_id_MPORT_mask = 1'h1;
  assign ram_class_meta_field_type_20_sub_class_id_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_class_meta_field_type_21_is_repeated_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_class_meta_field_type_21_is_repeated_io_deq_bits_MPORT_data =
    ram_class_meta_field_type_21_is_repeated[ram_class_meta_field_type_21_is_repeated_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  assign ram_class_meta_field_type_21_is_repeated_MPORT_data = io_enq_bits_class_meta_field_type_21_is_repeated;
  assign ram_class_meta_field_type_21_is_repeated_MPORT_addr = enq_ptr_value;
  assign ram_class_meta_field_type_21_is_repeated_MPORT_mask = 1'h1;
  assign ram_class_meta_field_type_21_is_repeated_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_class_meta_field_type_21_field_type_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_class_meta_field_type_21_field_type_io_deq_bits_MPORT_data =
    ram_class_meta_field_type_21_field_type[ram_class_meta_field_type_21_field_type_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  assign ram_class_meta_field_type_21_field_type_MPORT_data = io_enq_bits_class_meta_field_type_21_field_type;
  assign ram_class_meta_field_type_21_field_type_MPORT_addr = enq_ptr_value;
  assign ram_class_meta_field_type_21_field_type_MPORT_mask = 1'h1;
  assign ram_class_meta_field_type_21_field_type_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_class_meta_field_type_21_sub_class_id_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_class_meta_field_type_21_sub_class_id_io_deq_bits_MPORT_data =
    ram_class_meta_field_type_21_sub_class_id[ram_class_meta_field_type_21_sub_class_id_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  assign ram_class_meta_field_type_21_sub_class_id_MPORT_data = io_enq_bits_class_meta_field_type_21_sub_class_id;
  assign ram_class_meta_field_type_21_sub_class_id_MPORT_addr = enq_ptr_value;
  assign ram_class_meta_field_type_21_sub_class_id_MPORT_mask = 1'h1;
  assign ram_class_meta_field_type_21_sub_class_id_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_class_meta_field_type_22_is_repeated_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_class_meta_field_type_22_is_repeated_io_deq_bits_MPORT_data =
    ram_class_meta_field_type_22_is_repeated[ram_class_meta_field_type_22_is_repeated_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  assign ram_class_meta_field_type_22_is_repeated_MPORT_data = io_enq_bits_class_meta_field_type_22_is_repeated;
  assign ram_class_meta_field_type_22_is_repeated_MPORT_addr = enq_ptr_value;
  assign ram_class_meta_field_type_22_is_repeated_MPORT_mask = 1'h1;
  assign ram_class_meta_field_type_22_is_repeated_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_class_meta_field_type_22_field_type_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_class_meta_field_type_22_field_type_io_deq_bits_MPORT_data =
    ram_class_meta_field_type_22_field_type[ram_class_meta_field_type_22_field_type_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  assign ram_class_meta_field_type_22_field_type_MPORT_data = io_enq_bits_class_meta_field_type_22_field_type;
  assign ram_class_meta_field_type_22_field_type_MPORT_addr = enq_ptr_value;
  assign ram_class_meta_field_type_22_field_type_MPORT_mask = 1'h1;
  assign ram_class_meta_field_type_22_field_type_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_class_meta_field_type_22_sub_class_id_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_class_meta_field_type_22_sub_class_id_io_deq_bits_MPORT_data =
    ram_class_meta_field_type_22_sub_class_id[ram_class_meta_field_type_22_sub_class_id_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  assign ram_class_meta_field_type_22_sub_class_id_MPORT_data = io_enq_bits_class_meta_field_type_22_sub_class_id;
  assign ram_class_meta_field_type_22_sub_class_id_MPORT_addr = enq_ptr_value;
  assign ram_class_meta_field_type_22_sub_class_id_MPORT_mask = 1'h1;
  assign ram_class_meta_field_type_22_sub_class_id_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_class_meta_field_type_23_is_repeated_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_class_meta_field_type_23_is_repeated_io_deq_bits_MPORT_data =
    ram_class_meta_field_type_23_is_repeated[ram_class_meta_field_type_23_is_repeated_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  assign ram_class_meta_field_type_23_is_repeated_MPORT_data = io_enq_bits_class_meta_field_type_23_is_repeated;
  assign ram_class_meta_field_type_23_is_repeated_MPORT_addr = enq_ptr_value;
  assign ram_class_meta_field_type_23_is_repeated_MPORT_mask = 1'h1;
  assign ram_class_meta_field_type_23_is_repeated_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_class_meta_field_type_23_field_type_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_class_meta_field_type_23_field_type_io_deq_bits_MPORT_data =
    ram_class_meta_field_type_23_field_type[ram_class_meta_field_type_23_field_type_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  assign ram_class_meta_field_type_23_field_type_MPORT_data = io_enq_bits_class_meta_field_type_23_field_type;
  assign ram_class_meta_field_type_23_field_type_MPORT_addr = enq_ptr_value;
  assign ram_class_meta_field_type_23_field_type_MPORT_mask = 1'h1;
  assign ram_class_meta_field_type_23_field_type_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_class_meta_field_type_23_sub_class_id_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_class_meta_field_type_23_sub_class_id_io_deq_bits_MPORT_data =
    ram_class_meta_field_type_23_sub_class_id[ram_class_meta_field_type_23_sub_class_id_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  assign ram_class_meta_field_type_23_sub_class_id_MPORT_data = io_enq_bits_class_meta_field_type_23_sub_class_id;
  assign ram_class_meta_field_type_23_sub_class_id_MPORT_addr = enq_ptr_value;
  assign ram_class_meta_field_type_23_sub_class_id_MPORT_mask = 1'h1;
  assign ram_class_meta_field_type_23_sub_class_id_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_class_meta_field_type_24_is_repeated_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_class_meta_field_type_24_is_repeated_io_deq_bits_MPORT_data =
    ram_class_meta_field_type_24_is_repeated[ram_class_meta_field_type_24_is_repeated_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  assign ram_class_meta_field_type_24_is_repeated_MPORT_data = io_enq_bits_class_meta_field_type_24_is_repeated;
  assign ram_class_meta_field_type_24_is_repeated_MPORT_addr = enq_ptr_value;
  assign ram_class_meta_field_type_24_is_repeated_MPORT_mask = 1'h1;
  assign ram_class_meta_field_type_24_is_repeated_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_class_meta_field_type_24_field_type_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_class_meta_field_type_24_field_type_io_deq_bits_MPORT_data =
    ram_class_meta_field_type_24_field_type[ram_class_meta_field_type_24_field_type_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  assign ram_class_meta_field_type_24_field_type_MPORT_data = io_enq_bits_class_meta_field_type_24_field_type;
  assign ram_class_meta_field_type_24_field_type_MPORT_addr = enq_ptr_value;
  assign ram_class_meta_field_type_24_field_type_MPORT_mask = 1'h1;
  assign ram_class_meta_field_type_24_field_type_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_class_meta_field_type_24_sub_class_id_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_class_meta_field_type_24_sub_class_id_io_deq_bits_MPORT_data =
    ram_class_meta_field_type_24_sub_class_id[ram_class_meta_field_type_24_sub_class_id_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  assign ram_class_meta_field_type_24_sub_class_id_MPORT_data = io_enq_bits_class_meta_field_type_24_sub_class_id;
  assign ram_class_meta_field_type_24_sub_class_id_MPORT_addr = enq_ptr_value;
  assign ram_class_meta_field_type_24_sub_class_id_MPORT_mask = 1'h1;
  assign ram_class_meta_field_type_24_sub_class_id_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_class_meta_field_type_25_is_repeated_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_class_meta_field_type_25_is_repeated_io_deq_bits_MPORT_data =
    ram_class_meta_field_type_25_is_repeated[ram_class_meta_field_type_25_is_repeated_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  assign ram_class_meta_field_type_25_is_repeated_MPORT_data = io_enq_bits_class_meta_field_type_25_is_repeated;
  assign ram_class_meta_field_type_25_is_repeated_MPORT_addr = enq_ptr_value;
  assign ram_class_meta_field_type_25_is_repeated_MPORT_mask = 1'h1;
  assign ram_class_meta_field_type_25_is_repeated_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_class_meta_field_type_25_field_type_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_class_meta_field_type_25_field_type_io_deq_bits_MPORT_data =
    ram_class_meta_field_type_25_field_type[ram_class_meta_field_type_25_field_type_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  assign ram_class_meta_field_type_25_field_type_MPORT_data = io_enq_bits_class_meta_field_type_25_field_type;
  assign ram_class_meta_field_type_25_field_type_MPORT_addr = enq_ptr_value;
  assign ram_class_meta_field_type_25_field_type_MPORT_mask = 1'h1;
  assign ram_class_meta_field_type_25_field_type_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_class_meta_field_type_25_sub_class_id_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_class_meta_field_type_25_sub_class_id_io_deq_bits_MPORT_data =
    ram_class_meta_field_type_25_sub_class_id[ram_class_meta_field_type_25_sub_class_id_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  assign ram_class_meta_field_type_25_sub_class_id_MPORT_data = io_enq_bits_class_meta_field_type_25_sub_class_id;
  assign ram_class_meta_field_type_25_sub_class_id_MPORT_addr = enq_ptr_value;
  assign ram_class_meta_field_type_25_sub_class_id_MPORT_mask = 1'h1;
  assign ram_class_meta_field_type_25_sub_class_id_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_class_meta_field_type_26_is_repeated_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_class_meta_field_type_26_is_repeated_io_deq_bits_MPORT_data =
    ram_class_meta_field_type_26_is_repeated[ram_class_meta_field_type_26_is_repeated_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  assign ram_class_meta_field_type_26_is_repeated_MPORT_data = io_enq_bits_class_meta_field_type_26_is_repeated;
  assign ram_class_meta_field_type_26_is_repeated_MPORT_addr = enq_ptr_value;
  assign ram_class_meta_field_type_26_is_repeated_MPORT_mask = 1'h1;
  assign ram_class_meta_field_type_26_is_repeated_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_class_meta_field_type_26_field_type_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_class_meta_field_type_26_field_type_io_deq_bits_MPORT_data =
    ram_class_meta_field_type_26_field_type[ram_class_meta_field_type_26_field_type_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  assign ram_class_meta_field_type_26_field_type_MPORT_data = io_enq_bits_class_meta_field_type_26_field_type;
  assign ram_class_meta_field_type_26_field_type_MPORT_addr = enq_ptr_value;
  assign ram_class_meta_field_type_26_field_type_MPORT_mask = 1'h1;
  assign ram_class_meta_field_type_26_field_type_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_class_meta_field_type_26_sub_class_id_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_class_meta_field_type_26_sub_class_id_io_deq_bits_MPORT_data =
    ram_class_meta_field_type_26_sub_class_id[ram_class_meta_field_type_26_sub_class_id_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  assign ram_class_meta_field_type_26_sub_class_id_MPORT_data = io_enq_bits_class_meta_field_type_26_sub_class_id;
  assign ram_class_meta_field_type_26_sub_class_id_MPORT_addr = enq_ptr_value;
  assign ram_class_meta_field_type_26_sub_class_id_MPORT_mask = 1'h1;
  assign ram_class_meta_field_type_26_sub_class_id_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_class_meta_field_type_27_is_repeated_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_class_meta_field_type_27_is_repeated_io_deq_bits_MPORT_data =
    ram_class_meta_field_type_27_is_repeated[ram_class_meta_field_type_27_is_repeated_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  assign ram_class_meta_field_type_27_is_repeated_MPORT_data = io_enq_bits_class_meta_field_type_27_is_repeated;
  assign ram_class_meta_field_type_27_is_repeated_MPORT_addr = enq_ptr_value;
  assign ram_class_meta_field_type_27_is_repeated_MPORT_mask = 1'h1;
  assign ram_class_meta_field_type_27_is_repeated_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_class_meta_field_type_27_field_type_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_class_meta_field_type_27_field_type_io_deq_bits_MPORT_data =
    ram_class_meta_field_type_27_field_type[ram_class_meta_field_type_27_field_type_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  assign ram_class_meta_field_type_27_field_type_MPORT_data = io_enq_bits_class_meta_field_type_27_field_type;
  assign ram_class_meta_field_type_27_field_type_MPORT_addr = enq_ptr_value;
  assign ram_class_meta_field_type_27_field_type_MPORT_mask = 1'h1;
  assign ram_class_meta_field_type_27_field_type_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_class_meta_field_type_27_sub_class_id_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_class_meta_field_type_27_sub_class_id_io_deq_bits_MPORT_data =
    ram_class_meta_field_type_27_sub_class_id[ram_class_meta_field_type_27_sub_class_id_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  assign ram_class_meta_field_type_27_sub_class_id_MPORT_data = io_enq_bits_class_meta_field_type_27_sub_class_id;
  assign ram_class_meta_field_type_27_sub_class_id_MPORT_addr = enq_ptr_value;
  assign ram_class_meta_field_type_27_sub_class_id_MPORT_mask = 1'h1;
  assign ram_class_meta_field_type_27_sub_class_id_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_class_meta_field_type_28_is_repeated_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_class_meta_field_type_28_is_repeated_io_deq_bits_MPORT_data =
    ram_class_meta_field_type_28_is_repeated[ram_class_meta_field_type_28_is_repeated_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  assign ram_class_meta_field_type_28_is_repeated_MPORT_data = io_enq_bits_class_meta_field_type_28_is_repeated;
  assign ram_class_meta_field_type_28_is_repeated_MPORT_addr = enq_ptr_value;
  assign ram_class_meta_field_type_28_is_repeated_MPORT_mask = 1'h1;
  assign ram_class_meta_field_type_28_is_repeated_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_class_meta_field_type_28_field_type_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_class_meta_field_type_28_field_type_io_deq_bits_MPORT_data =
    ram_class_meta_field_type_28_field_type[ram_class_meta_field_type_28_field_type_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  assign ram_class_meta_field_type_28_field_type_MPORT_data = io_enq_bits_class_meta_field_type_28_field_type;
  assign ram_class_meta_field_type_28_field_type_MPORT_addr = enq_ptr_value;
  assign ram_class_meta_field_type_28_field_type_MPORT_mask = 1'h1;
  assign ram_class_meta_field_type_28_field_type_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_class_meta_field_type_28_sub_class_id_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_class_meta_field_type_28_sub_class_id_io_deq_bits_MPORT_data =
    ram_class_meta_field_type_28_sub_class_id[ram_class_meta_field_type_28_sub_class_id_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  assign ram_class_meta_field_type_28_sub_class_id_MPORT_data = io_enq_bits_class_meta_field_type_28_sub_class_id;
  assign ram_class_meta_field_type_28_sub_class_id_MPORT_addr = enq_ptr_value;
  assign ram_class_meta_field_type_28_sub_class_id_MPORT_mask = 1'h1;
  assign ram_class_meta_field_type_28_sub_class_id_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_class_meta_field_type_29_is_repeated_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_class_meta_field_type_29_is_repeated_io_deq_bits_MPORT_data =
    ram_class_meta_field_type_29_is_repeated[ram_class_meta_field_type_29_is_repeated_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  assign ram_class_meta_field_type_29_is_repeated_MPORT_data = io_enq_bits_class_meta_field_type_29_is_repeated;
  assign ram_class_meta_field_type_29_is_repeated_MPORT_addr = enq_ptr_value;
  assign ram_class_meta_field_type_29_is_repeated_MPORT_mask = 1'h1;
  assign ram_class_meta_field_type_29_is_repeated_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_class_meta_field_type_29_field_type_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_class_meta_field_type_29_field_type_io_deq_bits_MPORT_data =
    ram_class_meta_field_type_29_field_type[ram_class_meta_field_type_29_field_type_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  assign ram_class_meta_field_type_29_field_type_MPORT_data = io_enq_bits_class_meta_field_type_29_field_type;
  assign ram_class_meta_field_type_29_field_type_MPORT_addr = enq_ptr_value;
  assign ram_class_meta_field_type_29_field_type_MPORT_mask = 1'h1;
  assign ram_class_meta_field_type_29_field_type_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_class_meta_field_type_29_sub_class_id_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_class_meta_field_type_29_sub_class_id_io_deq_bits_MPORT_data =
    ram_class_meta_field_type_29_sub_class_id[ram_class_meta_field_type_29_sub_class_id_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  assign ram_class_meta_field_type_29_sub_class_id_MPORT_data = io_enq_bits_class_meta_field_type_29_sub_class_id;
  assign ram_class_meta_field_type_29_sub_class_id_MPORT_addr = enq_ptr_value;
  assign ram_class_meta_field_type_29_sub_class_id_MPORT_mask = 1'h1;
  assign ram_class_meta_field_type_29_sub_class_id_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_class_meta_field_type_30_is_repeated_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_class_meta_field_type_30_is_repeated_io_deq_bits_MPORT_data =
    ram_class_meta_field_type_30_is_repeated[ram_class_meta_field_type_30_is_repeated_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  assign ram_class_meta_field_type_30_is_repeated_MPORT_data = io_enq_bits_class_meta_field_type_30_is_repeated;
  assign ram_class_meta_field_type_30_is_repeated_MPORT_addr = enq_ptr_value;
  assign ram_class_meta_field_type_30_is_repeated_MPORT_mask = 1'h1;
  assign ram_class_meta_field_type_30_is_repeated_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_class_meta_field_type_30_field_type_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_class_meta_field_type_30_field_type_io_deq_bits_MPORT_data =
    ram_class_meta_field_type_30_field_type[ram_class_meta_field_type_30_field_type_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  assign ram_class_meta_field_type_30_field_type_MPORT_data = io_enq_bits_class_meta_field_type_30_field_type;
  assign ram_class_meta_field_type_30_field_type_MPORT_addr = enq_ptr_value;
  assign ram_class_meta_field_type_30_field_type_MPORT_mask = 1'h1;
  assign ram_class_meta_field_type_30_field_type_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_class_meta_field_type_30_sub_class_id_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_class_meta_field_type_30_sub_class_id_io_deq_bits_MPORT_data =
    ram_class_meta_field_type_30_sub_class_id[ram_class_meta_field_type_30_sub_class_id_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  assign ram_class_meta_field_type_30_sub_class_id_MPORT_data = io_enq_bits_class_meta_field_type_30_sub_class_id;
  assign ram_class_meta_field_type_30_sub_class_id_MPORT_addr = enq_ptr_value;
  assign ram_class_meta_field_type_30_sub_class_id_MPORT_mask = 1'h1;
  assign ram_class_meta_field_type_30_sub_class_id_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_class_meta_field_type_31_is_repeated_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_class_meta_field_type_31_is_repeated_io_deq_bits_MPORT_data =
    ram_class_meta_field_type_31_is_repeated[ram_class_meta_field_type_31_is_repeated_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  assign ram_class_meta_field_type_31_is_repeated_MPORT_data = io_enq_bits_class_meta_field_type_31_is_repeated;
  assign ram_class_meta_field_type_31_is_repeated_MPORT_addr = enq_ptr_value;
  assign ram_class_meta_field_type_31_is_repeated_MPORT_mask = 1'h1;
  assign ram_class_meta_field_type_31_is_repeated_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_class_meta_field_type_31_field_type_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_class_meta_field_type_31_field_type_io_deq_bits_MPORT_data =
    ram_class_meta_field_type_31_field_type[ram_class_meta_field_type_31_field_type_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  assign ram_class_meta_field_type_31_field_type_MPORT_data = io_enq_bits_class_meta_field_type_31_field_type;
  assign ram_class_meta_field_type_31_field_type_MPORT_addr = enq_ptr_value;
  assign ram_class_meta_field_type_31_field_type_MPORT_mask = 1'h1;
  assign ram_class_meta_field_type_31_field_type_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_class_meta_field_type_31_sub_class_id_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_class_meta_field_type_31_sub_class_id_io_deq_bits_MPORT_data =
    ram_class_meta_field_type_31_sub_class_id[ram_class_meta_field_type_31_sub_class_id_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  assign ram_class_meta_field_type_31_sub_class_id_MPORT_data = io_enq_bits_class_meta_field_type_31_sub_class_id;
  assign ram_class_meta_field_type_31_sub_class_id_MPORT_addr = enq_ptr_value;
  assign ram_class_meta_field_type_31_sub_class_id_MPORT_mask = 1'h1;
  assign ram_class_meta_field_type_31_sub_class_id_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_class_meta_field_type_32_is_repeated_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_class_meta_field_type_32_is_repeated_io_deq_bits_MPORT_data =
    ram_class_meta_field_type_32_is_repeated[ram_class_meta_field_type_32_is_repeated_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  assign ram_class_meta_field_type_32_is_repeated_MPORT_data = io_enq_bits_class_meta_field_type_32_is_repeated;
  assign ram_class_meta_field_type_32_is_repeated_MPORT_addr = enq_ptr_value;
  assign ram_class_meta_field_type_32_is_repeated_MPORT_mask = 1'h1;
  assign ram_class_meta_field_type_32_is_repeated_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_class_meta_field_type_32_field_type_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_class_meta_field_type_32_field_type_io_deq_bits_MPORT_data =
    ram_class_meta_field_type_32_field_type[ram_class_meta_field_type_32_field_type_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  assign ram_class_meta_field_type_32_field_type_MPORT_data = io_enq_bits_class_meta_field_type_32_field_type;
  assign ram_class_meta_field_type_32_field_type_MPORT_addr = enq_ptr_value;
  assign ram_class_meta_field_type_32_field_type_MPORT_mask = 1'h1;
  assign ram_class_meta_field_type_32_field_type_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_class_meta_field_type_32_sub_class_id_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_class_meta_field_type_32_sub_class_id_io_deq_bits_MPORT_data =
    ram_class_meta_field_type_32_sub_class_id[ram_class_meta_field_type_32_sub_class_id_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  assign ram_class_meta_field_type_32_sub_class_id_MPORT_data = io_enq_bits_class_meta_field_type_32_sub_class_id;
  assign ram_class_meta_field_type_32_sub_class_id_MPORT_addr = enq_ptr_value;
  assign ram_class_meta_field_type_32_sub_class_id_MPORT_mask = 1'h1;
  assign ram_class_meta_field_type_32_sub_class_id_MPORT_en = io_enq_ready & io_enq_valid;
  assign io_enq_ready = ~full; // @[Decoupled.scala 241:19]
  assign io_deq_valid = ~empty; // @[Decoupled.scala 240:19]
  assign io_deq_bits_class_meta_max_field_num = ram_class_meta_max_field_num_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15]
  assign io_deq_bits_class_meta_field_type_0_is_repeated =
    ram_class_meta_field_type_0_is_repeated_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15]
  assign io_deq_bits_class_meta_field_type_0_field_type = ram_class_meta_field_type_0_field_type_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15]
  assign io_deq_bits_class_meta_field_type_0_sub_class_id =
    ram_class_meta_field_type_0_sub_class_id_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15]
  assign io_deq_bits_class_meta_field_type_1_is_repeated =
    ram_class_meta_field_type_1_is_repeated_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15]
  assign io_deq_bits_class_meta_field_type_1_field_type = ram_class_meta_field_type_1_field_type_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15]
  assign io_deq_bits_class_meta_field_type_1_sub_class_id =
    ram_class_meta_field_type_1_sub_class_id_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15]
  assign io_deq_bits_class_meta_field_type_2_is_repeated =
    ram_class_meta_field_type_2_is_repeated_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15]
  assign io_deq_bits_class_meta_field_type_2_field_type = ram_class_meta_field_type_2_field_type_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15]
  assign io_deq_bits_class_meta_field_type_2_sub_class_id =
    ram_class_meta_field_type_2_sub_class_id_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15]
  assign io_deq_bits_class_meta_field_type_3_is_repeated =
    ram_class_meta_field_type_3_is_repeated_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15]
  assign io_deq_bits_class_meta_field_type_3_field_type = ram_class_meta_field_type_3_field_type_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15]
  assign io_deq_bits_class_meta_field_type_3_sub_class_id =
    ram_class_meta_field_type_3_sub_class_id_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15]
  assign io_deq_bits_class_meta_field_type_4_is_repeated =
    ram_class_meta_field_type_4_is_repeated_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15]
  assign io_deq_bits_class_meta_field_type_4_field_type = ram_class_meta_field_type_4_field_type_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15]
  assign io_deq_bits_class_meta_field_type_4_sub_class_id =
    ram_class_meta_field_type_4_sub_class_id_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15]
  assign io_deq_bits_class_meta_field_type_5_is_repeated =
    ram_class_meta_field_type_5_is_repeated_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15]
  assign io_deq_bits_class_meta_field_type_5_field_type = ram_class_meta_field_type_5_field_type_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15]
  assign io_deq_bits_class_meta_field_type_5_sub_class_id =
    ram_class_meta_field_type_5_sub_class_id_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15]
  assign io_deq_bits_class_meta_field_type_6_is_repeated =
    ram_class_meta_field_type_6_is_repeated_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15]
  assign io_deq_bits_class_meta_field_type_6_field_type = ram_class_meta_field_type_6_field_type_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15]
  assign io_deq_bits_class_meta_field_type_6_sub_class_id =
    ram_class_meta_field_type_6_sub_class_id_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15]
  assign io_deq_bits_class_meta_field_type_7_is_repeated =
    ram_class_meta_field_type_7_is_repeated_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15]
  assign io_deq_bits_class_meta_field_type_7_field_type = ram_class_meta_field_type_7_field_type_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15]
  assign io_deq_bits_class_meta_field_type_7_sub_class_id =
    ram_class_meta_field_type_7_sub_class_id_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15]
  assign io_deq_bits_class_meta_field_type_8_is_repeated =
    ram_class_meta_field_type_8_is_repeated_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15]
  assign io_deq_bits_class_meta_field_type_8_field_type = ram_class_meta_field_type_8_field_type_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15]
  assign io_deq_bits_class_meta_field_type_8_sub_class_id =
    ram_class_meta_field_type_8_sub_class_id_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15]
  assign io_deq_bits_class_meta_field_type_9_is_repeated =
    ram_class_meta_field_type_9_is_repeated_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15]
  assign io_deq_bits_class_meta_field_type_9_field_type = ram_class_meta_field_type_9_field_type_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15]
  assign io_deq_bits_class_meta_field_type_9_sub_class_id =
    ram_class_meta_field_type_9_sub_class_id_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15]
  assign io_deq_bits_class_meta_field_type_10_is_repeated =
    ram_class_meta_field_type_10_is_repeated_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15]
  assign io_deq_bits_class_meta_field_type_10_field_type =
    ram_class_meta_field_type_10_field_type_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15]
  assign io_deq_bits_class_meta_field_type_10_sub_class_id =
    ram_class_meta_field_type_10_sub_class_id_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15]
  assign io_deq_bits_class_meta_field_type_11_is_repeated =
    ram_class_meta_field_type_11_is_repeated_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15]
  assign io_deq_bits_class_meta_field_type_11_field_type =
    ram_class_meta_field_type_11_field_type_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15]
  assign io_deq_bits_class_meta_field_type_11_sub_class_id =
    ram_class_meta_field_type_11_sub_class_id_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15]
  assign io_deq_bits_class_meta_field_type_12_is_repeated =
    ram_class_meta_field_type_12_is_repeated_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15]
  assign io_deq_bits_class_meta_field_type_12_field_type =
    ram_class_meta_field_type_12_field_type_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15]
  assign io_deq_bits_class_meta_field_type_12_sub_class_id =
    ram_class_meta_field_type_12_sub_class_id_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15]
  assign io_deq_bits_class_meta_field_type_13_is_repeated =
    ram_class_meta_field_type_13_is_repeated_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15]
  assign io_deq_bits_class_meta_field_type_13_field_type =
    ram_class_meta_field_type_13_field_type_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15]
  assign io_deq_bits_class_meta_field_type_13_sub_class_id =
    ram_class_meta_field_type_13_sub_class_id_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15]
  assign io_deq_bits_class_meta_field_type_14_is_repeated =
    ram_class_meta_field_type_14_is_repeated_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15]
  assign io_deq_bits_class_meta_field_type_14_field_type =
    ram_class_meta_field_type_14_field_type_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15]
  assign io_deq_bits_class_meta_field_type_14_sub_class_id =
    ram_class_meta_field_type_14_sub_class_id_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15]
  assign io_deq_bits_class_meta_field_type_15_is_repeated =
    ram_class_meta_field_type_15_is_repeated_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15]
  assign io_deq_bits_class_meta_field_type_15_field_type =
    ram_class_meta_field_type_15_field_type_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15]
  assign io_deq_bits_class_meta_field_type_15_sub_class_id =
    ram_class_meta_field_type_15_sub_class_id_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15]
  assign io_deq_bits_class_meta_field_type_16_is_repeated =
    ram_class_meta_field_type_16_is_repeated_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15]
  assign io_deq_bits_class_meta_field_type_16_field_type =
    ram_class_meta_field_type_16_field_type_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15]
  assign io_deq_bits_class_meta_field_type_16_sub_class_id =
    ram_class_meta_field_type_16_sub_class_id_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15]
  assign io_deq_bits_class_meta_field_type_17_is_repeated =
    ram_class_meta_field_type_17_is_repeated_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15]
  assign io_deq_bits_class_meta_field_type_17_field_type =
    ram_class_meta_field_type_17_field_type_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15]
  assign io_deq_bits_class_meta_field_type_17_sub_class_id =
    ram_class_meta_field_type_17_sub_class_id_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15]
  assign io_deq_bits_class_meta_field_type_18_is_repeated =
    ram_class_meta_field_type_18_is_repeated_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15]
  assign io_deq_bits_class_meta_field_type_18_field_type =
    ram_class_meta_field_type_18_field_type_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15]
  assign io_deq_bits_class_meta_field_type_18_sub_class_id =
    ram_class_meta_field_type_18_sub_class_id_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15]
  assign io_deq_bits_class_meta_field_type_19_is_repeated =
    ram_class_meta_field_type_19_is_repeated_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15]
  assign io_deq_bits_class_meta_field_type_19_field_type =
    ram_class_meta_field_type_19_field_type_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15]
  assign io_deq_bits_class_meta_field_type_19_sub_class_id =
    ram_class_meta_field_type_19_sub_class_id_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15]
  assign io_deq_bits_class_meta_field_type_20_is_repeated =
    ram_class_meta_field_type_20_is_repeated_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15]
  assign io_deq_bits_class_meta_field_type_20_field_type =
    ram_class_meta_field_type_20_field_type_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15]
  assign io_deq_bits_class_meta_field_type_20_sub_class_id =
    ram_class_meta_field_type_20_sub_class_id_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15]
  assign io_deq_bits_class_meta_field_type_21_is_repeated =
    ram_class_meta_field_type_21_is_repeated_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15]
  assign io_deq_bits_class_meta_field_type_21_field_type =
    ram_class_meta_field_type_21_field_type_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15]
  assign io_deq_bits_class_meta_field_type_21_sub_class_id =
    ram_class_meta_field_type_21_sub_class_id_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15]
  assign io_deq_bits_class_meta_field_type_22_is_repeated =
    ram_class_meta_field_type_22_is_repeated_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15]
  assign io_deq_bits_class_meta_field_type_22_field_type =
    ram_class_meta_field_type_22_field_type_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15]
  assign io_deq_bits_class_meta_field_type_22_sub_class_id =
    ram_class_meta_field_type_22_sub_class_id_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15]
  assign io_deq_bits_class_meta_field_type_23_is_repeated =
    ram_class_meta_field_type_23_is_repeated_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15]
  assign io_deq_bits_class_meta_field_type_23_field_type =
    ram_class_meta_field_type_23_field_type_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15]
  assign io_deq_bits_class_meta_field_type_23_sub_class_id =
    ram_class_meta_field_type_23_sub_class_id_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15]
  assign io_deq_bits_class_meta_field_type_24_is_repeated =
    ram_class_meta_field_type_24_is_repeated_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15]
  assign io_deq_bits_class_meta_field_type_24_field_type =
    ram_class_meta_field_type_24_field_type_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15]
  assign io_deq_bits_class_meta_field_type_24_sub_class_id =
    ram_class_meta_field_type_24_sub_class_id_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15]
  assign io_deq_bits_class_meta_field_type_25_is_repeated =
    ram_class_meta_field_type_25_is_repeated_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15]
  assign io_deq_bits_class_meta_field_type_25_field_type =
    ram_class_meta_field_type_25_field_type_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15]
  assign io_deq_bits_class_meta_field_type_25_sub_class_id =
    ram_class_meta_field_type_25_sub_class_id_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15]
  assign io_deq_bits_class_meta_field_type_26_is_repeated =
    ram_class_meta_field_type_26_is_repeated_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15]
  assign io_deq_bits_class_meta_field_type_26_field_type =
    ram_class_meta_field_type_26_field_type_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15]
  assign io_deq_bits_class_meta_field_type_26_sub_class_id =
    ram_class_meta_field_type_26_sub_class_id_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15]
  assign io_deq_bits_class_meta_field_type_27_is_repeated =
    ram_class_meta_field_type_27_is_repeated_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15]
  assign io_deq_bits_class_meta_field_type_27_field_type =
    ram_class_meta_field_type_27_field_type_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15]
  assign io_deq_bits_class_meta_field_type_27_sub_class_id =
    ram_class_meta_field_type_27_sub_class_id_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15]
  assign io_deq_bits_class_meta_field_type_28_is_repeated =
    ram_class_meta_field_type_28_is_repeated_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15]
  assign io_deq_bits_class_meta_field_type_28_field_type =
    ram_class_meta_field_type_28_field_type_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15]
  assign io_deq_bits_class_meta_field_type_28_sub_class_id =
    ram_class_meta_field_type_28_sub_class_id_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15]
  assign io_deq_bits_class_meta_field_type_29_is_repeated =
    ram_class_meta_field_type_29_is_repeated_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15]
  assign io_deq_bits_class_meta_field_type_29_field_type =
    ram_class_meta_field_type_29_field_type_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15]
  assign io_deq_bits_class_meta_field_type_29_sub_class_id =
    ram_class_meta_field_type_29_sub_class_id_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15]
  assign io_deq_bits_class_meta_field_type_30_is_repeated =
    ram_class_meta_field_type_30_is_repeated_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15]
  assign io_deq_bits_class_meta_field_type_30_field_type =
    ram_class_meta_field_type_30_field_type_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15]
  assign io_deq_bits_class_meta_field_type_30_sub_class_id =
    ram_class_meta_field_type_30_sub_class_id_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15]
  assign io_deq_bits_class_meta_field_type_31_is_repeated =
    ram_class_meta_field_type_31_is_repeated_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15]
  assign io_deq_bits_class_meta_field_type_31_field_type =
    ram_class_meta_field_type_31_field_type_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15]
  assign io_deq_bits_class_meta_field_type_31_sub_class_id =
    ram_class_meta_field_type_31_sub_class_id_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15]
  assign io_deq_bits_class_meta_field_type_32_is_repeated =
    ram_class_meta_field_type_32_is_repeated_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15]
  assign io_deq_bits_class_meta_field_type_32_field_type =
    ram_class_meta_field_type_32_field_type_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15]
  assign io_deq_bits_class_meta_field_type_32_sub_class_id =
    ram_class_meta_field_type_32_sub_class_id_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15]
  always @(posedge clock) begin
    if(ram_class_meta_max_field_num_MPORT_en & ram_class_meta_max_field_num_MPORT_mask) begin
      ram_class_meta_max_field_num[ram_class_meta_max_field_num_MPORT_addr] <= ram_class_meta_max_field_num_MPORT_data; // @[Decoupled.scala 218:16]
    end
    if(ram_class_meta_field_type_0_is_repeated_MPORT_en & ram_class_meta_field_type_0_is_repeated_MPORT_mask) begin
      ram_class_meta_field_type_0_is_repeated[ram_class_meta_field_type_0_is_repeated_MPORT_addr] <=
        ram_class_meta_field_type_0_is_repeated_MPORT_data; // @[Decoupled.scala 218:16]
    end
    if(ram_class_meta_field_type_0_field_type_MPORT_en & ram_class_meta_field_type_0_field_type_MPORT_mask) begin
      ram_class_meta_field_type_0_field_type[ram_class_meta_field_type_0_field_type_MPORT_addr] <=
        ram_class_meta_field_type_0_field_type_MPORT_data; // @[Decoupled.scala 218:16]
    end
    if(ram_class_meta_field_type_0_sub_class_id_MPORT_en & ram_class_meta_field_type_0_sub_class_id_MPORT_mask) begin
      ram_class_meta_field_type_0_sub_class_id[ram_class_meta_field_type_0_sub_class_id_MPORT_addr] <=
        ram_class_meta_field_type_0_sub_class_id_MPORT_data; // @[Decoupled.scala 218:16]
    end
    if(ram_class_meta_field_type_1_is_repeated_MPORT_en & ram_class_meta_field_type_1_is_repeated_MPORT_mask) begin
      ram_class_meta_field_type_1_is_repeated[ram_class_meta_field_type_1_is_repeated_MPORT_addr] <=
        ram_class_meta_field_type_1_is_repeated_MPORT_data; // @[Decoupled.scala 218:16]
    end
    if(ram_class_meta_field_type_1_field_type_MPORT_en & ram_class_meta_field_type_1_field_type_MPORT_mask) begin
      ram_class_meta_field_type_1_field_type[ram_class_meta_field_type_1_field_type_MPORT_addr] <=
        ram_class_meta_field_type_1_field_type_MPORT_data; // @[Decoupled.scala 218:16]
    end
    if(ram_class_meta_field_type_1_sub_class_id_MPORT_en & ram_class_meta_field_type_1_sub_class_id_MPORT_mask) begin
      ram_class_meta_field_type_1_sub_class_id[ram_class_meta_field_type_1_sub_class_id_MPORT_addr] <=
        ram_class_meta_field_type_1_sub_class_id_MPORT_data; // @[Decoupled.scala 218:16]
    end
    if(ram_class_meta_field_type_2_is_repeated_MPORT_en & ram_class_meta_field_type_2_is_repeated_MPORT_mask) begin
      ram_class_meta_field_type_2_is_repeated[ram_class_meta_field_type_2_is_repeated_MPORT_addr] <=
        ram_class_meta_field_type_2_is_repeated_MPORT_data; // @[Decoupled.scala 218:16]
    end
    if(ram_class_meta_field_type_2_field_type_MPORT_en & ram_class_meta_field_type_2_field_type_MPORT_mask) begin
      ram_class_meta_field_type_2_field_type[ram_class_meta_field_type_2_field_type_MPORT_addr] <=
        ram_class_meta_field_type_2_field_type_MPORT_data; // @[Decoupled.scala 218:16]
    end
    if(ram_class_meta_field_type_2_sub_class_id_MPORT_en & ram_class_meta_field_type_2_sub_class_id_MPORT_mask) begin
      ram_class_meta_field_type_2_sub_class_id[ram_class_meta_field_type_2_sub_class_id_MPORT_addr] <=
        ram_class_meta_field_type_2_sub_class_id_MPORT_data; // @[Decoupled.scala 218:16]
    end
    if(ram_class_meta_field_type_3_is_repeated_MPORT_en & ram_class_meta_field_type_3_is_repeated_MPORT_mask) begin
      ram_class_meta_field_type_3_is_repeated[ram_class_meta_field_type_3_is_repeated_MPORT_addr] <=
        ram_class_meta_field_type_3_is_repeated_MPORT_data; // @[Decoupled.scala 218:16]
    end
    if(ram_class_meta_field_type_3_field_type_MPORT_en & ram_class_meta_field_type_3_field_type_MPORT_mask) begin
      ram_class_meta_field_type_3_field_type[ram_class_meta_field_type_3_field_type_MPORT_addr] <=
        ram_class_meta_field_type_3_field_type_MPORT_data; // @[Decoupled.scala 218:16]
    end
    if(ram_class_meta_field_type_3_sub_class_id_MPORT_en & ram_class_meta_field_type_3_sub_class_id_MPORT_mask) begin
      ram_class_meta_field_type_3_sub_class_id[ram_class_meta_field_type_3_sub_class_id_MPORT_addr] <=
        ram_class_meta_field_type_3_sub_class_id_MPORT_data; // @[Decoupled.scala 218:16]
    end
    if(ram_class_meta_field_type_4_is_repeated_MPORT_en & ram_class_meta_field_type_4_is_repeated_MPORT_mask) begin
      ram_class_meta_field_type_4_is_repeated[ram_class_meta_field_type_4_is_repeated_MPORT_addr] <=
        ram_class_meta_field_type_4_is_repeated_MPORT_data; // @[Decoupled.scala 218:16]
    end
    if(ram_class_meta_field_type_4_field_type_MPORT_en & ram_class_meta_field_type_4_field_type_MPORT_mask) begin
      ram_class_meta_field_type_4_field_type[ram_class_meta_field_type_4_field_type_MPORT_addr] <=
        ram_class_meta_field_type_4_field_type_MPORT_data; // @[Decoupled.scala 218:16]
    end
    if(ram_class_meta_field_type_4_sub_class_id_MPORT_en & ram_class_meta_field_type_4_sub_class_id_MPORT_mask) begin
      ram_class_meta_field_type_4_sub_class_id[ram_class_meta_field_type_4_sub_class_id_MPORT_addr] <=
        ram_class_meta_field_type_4_sub_class_id_MPORT_data; // @[Decoupled.scala 218:16]
    end
    if(ram_class_meta_field_type_5_is_repeated_MPORT_en & ram_class_meta_field_type_5_is_repeated_MPORT_mask) begin
      ram_class_meta_field_type_5_is_repeated[ram_class_meta_field_type_5_is_repeated_MPORT_addr] <=
        ram_class_meta_field_type_5_is_repeated_MPORT_data; // @[Decoupled.scala 218:16]
    end
    if(ram_class_meta_field_type_5_field_type_MPORT_en & ram_class_meta_field_type_5_field_type_MPORT_mask) begin
      ram_class_meta_field_type_5_field_type[ram_class_meta_field_type_5_field_type_MPORT_addr] <=
        ram_class_meta_field_type_5_field_type_MPORT_data; // @[Decoupled.scala 218:16]
    end
    if(ram_class_meta_field_type_5_sub_class_id_MPORT_en & ram_class_meta_field_type_5_sub_class_id_MPORT_mask) begin
      ram_class_meta_field_type_5_sub_class_id[ram_class_meta_field_type_5_sub_class_id_MPORT_addr] <=
        ram_class_meta_field_type_5_sub_class_id_MPORT_data; // @[Decoupled.scala 218:16]
    end
    if(ram_class_meta_field_type_6_is_repeated_MPORT_en & ram_class_meta_field_type_6_is_repeated_MPORT_mask) begin
      ram_class_meta_field_type_6_is_repeated[ram_class_meta_field_type_6_is_repeated_MPORT_addr] <=
        ram_class_meta_field_type_6_is_repeated_MPORT_data; // @[Decoupled.scala 218:16]
    end
    if(ram_class_meta_field_type_6_field_type_MPORT_en & ram_class_meta_field_type_6_field_type_MPORT_mask) begin
      ram_class_meta_field_type_6_field_type[ram_class_meta_field_type_6_field_type_MPORT_addr] <=
        ram_class_meta_field_type_6_field_type_MPORT_data; // @[Decoupled.scala 218:16]
    end
    if(ram_class_meta_field_type_6_sub_class_id_MPORT_en & ram_class_meta_field_type_6_sub_class_id_MPORT_mask) begin
      ram_class_meta_field_type_6_sub_class_id[ram_class_meta_field_type_6_sub_class_id_MPORT_addr] <=
        ram_class_meta_field_type_6_sub_class_id_MPORT_data; // @[Decoupled.scala 218:16]
    end
    if(ram_class_meta_field_type_7_is_repeated_MPORT_en & ram_class_meta_field_type_7_is_repeated_MPORT_mask) begin
      ram_class_meta_field_type_7_is_repeated[ram_class_meta_field_type_7_is_repeated_MPORT_addr] <=
        ram_class_meta_field_type_7_is_repeated_MPORT_data; // @[Decoupled.scala 218:16]
    end
    if(ram_class_meta_field_type_7_field_type_MPORT_en & ram_class_meta_field_type_7_field_type_MPORT_mask) begin
      ram_class_meta_field_type_7_field_type[ram_class_meta_field_type_7_field_type_MPORT_addr] <=
        ram_class_meta_field_type_7_field_type_MPORT_data; // @[Decoupled.scala 218:16]
    end
    if(ram_class_meta_field_type_7_sub_class_id_MPORT_en & ram_class_meta_field_type_7_sub_class_id_MPORT_mask) begin
      ram_class_meta_field_type_7_sub_class_id[ram_class_meta_field_type_7_sub_class_id_MPORT_addr] <=
        ram_class_meta_field_type_7_sub_class_id_MPORT_data; // @[Decoupled.scala 218:16]
    end
    if(ram_class_meta_field_type_8_is_repeated_MPORT_en & ram_class_meta_field_type_8_is_repeated_MPORT_mask) begin
      ram_class_meta_field_type_8_is_repeated[ram_class_meta_field_type_8_is_repeated_MPORT_addr] <=
        ram_class_meta_field_type_8_is_repeated_MPORT_data; // @[Decoupled.scala 218:16]
    end
    if(ram_class_meta_field_type_8_field_type_MPORT_en & ram_class_meta_field_type_8_field_type_MPORT_mask) begin
      ram_class_meta_field_type_8_field_type[ram_class_meta_field_type_8_field_type_MPORT_addr] <=
        ram_class_meta_field_type_8_field_type_MPORT_data; // @[Decoupled.scala 218:16]
    end
    if(ram_class_meta_field_type_8_sub_class_id_MPORT_en & ram_class_meta_field_type_8_sub_class_id_MPORT_mask) begin
      ram_class_meta_field_type_8_sub_class_id[ram_class_meta_field_type_8_sub_class_id_MPORT_addr] <=
        ram_class_meta_field_type_8_sub_class_id_MPORT_data; // @[Decoupled.scala 218:16]
    end
    if(ram_class_meta_field_type_9_is_repeated_MPORT_en & ram_class_meta_field_type_9_is_repeated_MPORT_mask) begin
      ram_class_meta_field_type_9_is_repeated[ram_class_meta_field_type_9_is_repeated_MPORT_addr] <=
        ram_class_meta_field_type_9_is_repeated_MPORT_data; // @[Decoupled.scala 218:16]
    end
    if(ram_class_meta_field_type_9_field_type_MPORT_en & ram_class_meta_field_type_9_field_type_MPORT_mask) begin
      ram_class_meta_field_type_9_field_type[ram_class_meta_field_type_9_field_type_MPORT_addr] <=
        ram_class_meta_field_type_9_field_type_MPORT_data; // @[Decoupled.scala 218:16]
    end
    if(ram_class_meta_field_type_9_sub_class_id_MPORT_en & ram_class_meta_field_type_9_sub_class_id_MPORT_mask) begin
      ram_class_meta_field_type_9_sub_class_id[ram_class_meta_field_type_9_sub_class_id_MPORT_addr] <=
        ram_class_meta_field_type_9_sub_class_id_MPORT_data; // @[Decoupled.scala 218:16]
    end
    if(ram_class_meta_field_type_10_is_repeated_MPORT_en & ram_class_meta_field_type_10_is_repeated_MPORT_mask) begin
      ram_class_meta_field_type_10_is_repeated[ram_class_meta_field_type_10_is_repeated_MPORT_addr] <=
        ram_class_meta_field_type_10_is_repeated_MPORT_data; // @[Decoupled.scala 218:16]
    end
    if(ram_class_meta_field_type_10_field_type_MPORT_en & ram_class_meta_field_type_10_field_type_MPORT_mask) begin
      ram_class_meta_field_type_10_field_type[ram_class_meta_field_type_10_field_type_MPORT_addr] <=
        ram_class_meta_field_type_10_field_type_MPORT_data; // @[Decoupled.scala 218:16]
    end
    if(ram_class_meta_field_type_10_sub_class_id_MPORT_en & ram_class_meta_field_type_10_sub_class_id_MPORT_mask) begin
      ram_class_meta_field_type_10_sub_class_id[ram_class_meta_field_type_10_sub_class_id_MPORT_addr] <=
        ram_class_meta_field_type_10_sub_class_id_MPORT_data; // @[Decoupled.scala 218:16]
    end
    if(ram_class_meta_field_type_11_is_repeated_MPORT_en & ram_class_meta_field_type_11_is_repeated_MPORT_mask) begin
      ram_class_meta_field_type_11_is_repeated[ram_class_meta_field_type_11_is_repeated_MPORT_addr] <=
        ram_class_meta_field_type_11_is_repeated_MPORT_data; // @[Decoupled.scala 218:16]
    end
    if(ram_class_meta_field_type_11_field_type_MPORT_en & ram_class_meta_field_type_11_field_type_MPORT_mask) begin
      ram_class_meta_field_type_11_field_type[ram_class_meta_field_type_11_field_type_MPORT_addr] <=
        ram_class_meta_field_type_11_field_type_MPORT_data; // @[Decoupled.scala 218:16]
    end
    if(ram_class_meta_field_type_11_sub_class_id_MPORT_en & ram_class_meta_field_type_11_sub_class_id_MPORT_mask) begin
      ram_class_meta_field_type_11_sub_class_id[ram_class_meta_field_type_11_sub_class_id_MPORT_addr] <=
        ram_class_meta_field_type_11_sub_class_id_MPORT_data; // @[Decoupled.scala 218:16]
    end
    if(ram_class_meta_field_type_12_is_repeated_MPORT_en & ram_class_meta_field_type_12_is_repeated_MPORT_mask) begin
      ram_class_meta_field_type_12_is_repeated[ram_class_meta_field_type_12_is_repeated_MPORT_addr] <=
        ram_class_meta_field_type_12_is_repeated_MPORT_data; // @[Decoupled.scala 218:16]
    end
    if(ram_class_meta_field_type_12_field_type_MPORT_en & ram_class_meta_field_type_12_field_type_MPORT_mask) begin
      ram_class_meta_field_type_12_field_type[ram_class_meta_field_type_12_field_type_MPORT_addr] <=
        ram_class_meta_field_type_12_field_type_MPORT_data; // @[Decoupled.scala 218:16]
    end
    if(ram_class_meta_field_type_12_sub_class_id_MPORT_en & ram_class_meta_field_type_12_sub_class_id_MPORT_mask) begin
      ram_class_meta_field_type_12_sub_class_id[ram_class_meta_field_type_12_sub_class_id_MPORT_addr] <=
        ram_class_meta_field_type_12_sub_class_id_MPORT_data; // @[Decoupled.scala 218:16]
    end
    if(ram_class_meta_field_type_13_is_repeated_MPORT_en & ram_class_meta_field_type_13_is_repeated_MPORT_mask) begin
      ram_class_meta_field_type_13_is_repeated[ram_class_meta_field_type_13_is_repeated_MPORT_addr] <=
        ram_class_meta_field_type_13_is_repeated_MPORT_data; // @[Decoupled.scala 218:16]
    end
    if(ram_class_meta_field_type_13_field_type_MPORT_en & ram_class_meta_field_type_13_field_type_MPORT_mask) begin
      ram_class_meta_field_type_13_field_type[ram_class_meta_field_type_13_field_type_MPORT_addr] <=
        ram_class_meta_field_type_13_field_type_MPORT_data; // @[Decoupled.scala 218:16]
    end
    if(ram_class_meta_field_type_13_sub_class_id_MPORT_en & ram_class_meta_field_type_13_sub_class_id_MPORT_mask) begin
      ram_class_meta_field_type_13_sub_class_id[ram_class_meta_field_type_13_sub_class_id_MPORT_addr] <=
        ram_class_meta_field_type_13_sub_class_id_MPORT_data; // @[Decoupled.scala 218:16]
    end
    if(ram_class_meta_field_type_14_is_repeated_MPORT_en & ram_class_meta_field_type_14_is_repeated_MPORT_mask) begin
      ram_class_meta_field_type_14_is_repeated[ram_class_meta_field_type_14_is_repeated_MPORT_addr] <=
        ram_class_meta_field_type_14_is_repeated_MPORT_data; // @[Decoupled.scala 218:16]
    end
    if(ram_class_meta_field_type_14_field_type_MPORT_en & ram_class_meta_field_type_14_field_type_MPORT_mask) begin
      ram_class_meta_field_type_14_field_type[ram_class_meta_field_type_14_field_type_MPORT_addr] <=
        ram_class_meta_field_type_14_field_type_MPORT_data; // @[Decoupled.scala 218:16]
    end
    if(ram_class_meta_field_type_14_sub_class_id_MPORT_en & ram_class_meta_field_type_14_sub_class_id_MPORT_mask) begin
      ram_class_meta_field_type_14_sub_class_id[ram_class_meta_field_type_14_sub_class_id_MPORT_addr] <=
        ram_class_meta_field_type_14_sub_class_id_MPORT_data; // @[Decoupled.scala 218:16]
    end
    if(ram_class_meta_field_type_15_is_repeated_MPORT_en & ram_class_meta_field_type_15_is_repeated_MPORT_mask) begin
      ram_class_meta_field_type_15_is_repeated[ram_class_meta_field_type_15_is_repeated_MPORT_addr] <=
        ram_class_meta_field_type_15_is_repeated_MPORT_data; // @[Decoupled.scala 218:16]
    end
    if(ram_class_meta_field_type_15_field_type_MPORT_en & ram_class_meta_field_type_15_field_type_MPORT_mask) begin
      ram_class_meta_field_type_15_field_type[ram_class_meta_field_type_15_field_type_MPORT_addr] <=
        ram_class_meta_field_type_15_field_type_MPORT_data; // @[Decoupled.scala 218:16]
    end
    if(ram_class_meta_field_type_15_sub_class_id_MPORT_en & ram_class_meta_field_type_15_sub_class_id_MPORT_mask) begin
      ram_class_meta_field_type_15_sub_class_id[ram_class_meta_field_type_15_sub_class_id_MPORT_addr] <=
        ram_class_meta_field_type_15_sub_class_id_MPORT_data; // @[Decoupled.scala 218:16]
    end
    if(ram_class_meta_field_type_16_is_repeated_MPORT_en & ram_class_meta_field_type_16_is_repeated_MPORT_mask) begin
      ram_class_meta_field_type_16_is_repeated[ram_class_meta_field_type_16_is_repeated_MPORT_addr] <=
        ram_class_meta_field_type_16_is_repeated_MPORT_data; // @[Decoupled.scala 218:16]
    end
    if(ram_class_meta_field_type_16_field_type_MPORT_en & ram_class_meta_field_type_16_field_type_MPORT_mask) begin
      ram_class_meta_field_type_16_field_type[ram_class_meta_field_type_16_field_type_MPORT_addr] <=
        ram_class_meta_field_type_16_field_type_MPORT_data; // @[Decoupled.scala 218:16]
    end
    if(ram_class_meta_field_type_16_sub_class_id_MPORT_en & ram_class_meta_field_type_16_sub_class_id_MPORT_mask) begin
      ram_class_meta_field_type_16_sub_class_id[ram_class_meta_field_type_16_sub_class_id_MPORT_addr] <=
        ram_class_meta_field_type_16_sub_class_id_MPORT_data; // @[Decoupled.scala 218:16]
    end
    if(ram_class_meta_field_type_17_is_repeated_MPORT_en & ram_class_meta_field_type_17_is_repeated_MPORT_mask) begin
      ram_class_meta_field_type_17_is_repeated[ram_class_meta_field_type_17_is_repeated_MPORT_addr] <=
        ram_class_meta_field_type_17_is_repeated_MPORT_data; // @[Decoupled.scala 218:16]
    end
    if(ram_class_meta_field_type_17_field_type_MPORT_en & ram_class_meta_field_type_17_field_type_MPORT_mask) begin
      ram_class_meta_field_type_17_field_type[ram_class_meta_field_type_17_field_type_MPORT_addr] <=
        ram_class_meta_field_type_17_field_type_MPORT_data; // @[Decoupled.scala 218:16]
    end
    if(ram_class_meta_field_type_17_sub_class_id_MPORT_en & ram_class_meta_field_type_17_sub_class_id_MPORT_mask) begin
      ram_class_meta_field_type_17_sub_class_id[ram_class_meta_field_type_17_sub_class_id_MPORT_addr] <=
        ram_class_meta_field_type_17_sub_class_id_MPORT_data; // @[Decoupled.scala 218:16]
    end
    if(ram_class_meta_field_type_18_is_repeated_MPORT_en & ram_class_meta_field_type_18_is_repeated_MPORT_mask) begin
      ram_class_meta_field_type_18_is_repeated[ram_class_meta_field_type_18_is_repeated_MPORT_addr] <=
        ram_class_meta_field_type_18_is_repeated_MPORT_data; // @[Decoupled.scala 218:16]
    end
    if(ram_class_meta_field_type_18_field_type_MPORT_en & ram_class_meta_field_type_18_field_type_MPORT_mask) begin
      ram_class_meta_field_type_18_field_type[ram_class_meta_field_type_18_field_type_MPORT_addr] <=
        ram_class_meta_field_type_18_field_type_MPORT_data; // @[Decoupled.scala 218:16]
    end
    if(ram_class_meta_field_type_18_sub_class_id_MPORT_en & ram_class_meta_field_type_18_sub_class_id_MPORT_mask) begin
      ram_class_meta_field_type_18_sub_class_id[ram_class_meta_field_type_18_sub_class_id_MPORT_addr] <=
        ram_class_meta_field_type_18_sub_class_id_MPORT_data; // @[Decoupled.scala 218:16]
    end
    if(ram_class_meta_field_type_19_is_repeated_MPORT_en & ram_class_meta_field_type_19_is_repeated_MPORT_mask) begin
      ram_class_meta_field_type_19_is_repeated[ram_class_meta_field_type_19_is_repeated_MPORT_addr] <=
        ram_class_meta_field_type_19_is_repeated_MPORT_data; // @[Decoupled.scala 218:16]
    end
    if(ram_class_meta_field_type_19_field_type_MPORT_en & ram_class_meta_field_type_19_field_type_MPORT_mask) begin
      ram_class_meta_field_type_19_field_type[ram_class_meta_field_type_19_field_type_MPORT_addr] <=
        ram_class_meta_field_type_19_field_type_MPORT_data; // @[Decoupled.scala 218:16]
    end
    if(ram_class_meta_field_type_19_sub_class_id_MPORT_en & ram_class_meta_field_type_19_sub_class_id_MPORT_mask) begin
      ram_class_meta_field_type_19_sub_class_id[ram_class_meta_field_type_19_sub_class_id_MPORT_addr] <=
        ram_class_meta_field_type_19_sub_class_id_MPORT_data; // @[Decoupled.scala 218:16]
    end
    if(ram_class_meta_field_type_20_is_repeated_MPORT_en & ram_class_meta_field_type_20_is_repeated_MPORT_mask) begin
      ram_class_meta_field_type_20_is_repeated[ram_class_meta_field_type_20_is_repeated_MPORT_addr] <=
        ram_class_meta_field_type_20_is_repeated_MPORT_data; // @[Decoupled.scala 218:16]
    end
    if(ram_class_meta_field_type_20_field_type_MPORT_en & ram_class_meta_field_type_20_field_type_MPORT_mask) begin
      ram_class_meta_field_type_20_field_type[ram_class_meta_field_type_20_field_type_MPORT_addr] <=
        ram_class_meta_field_type_20_field_type_MPORT_data; // @[Decoupled.scala 218:16]
    end
    if(ram_class_meta_field_type_20_sub_class_id_MPORT_en & ram_class_meta_field_type_20_sub_class_id_MPORT_mask) begin
      ram_class_meta_field_type_20_sub_class_id[ram_class_meta_field_type_20_sub_class_id_MPORT_addr] <=
        ram_class_meta_field_type_20_sub_class_id_MPORT_data; // @[Decoupled.scala 218:16]
    end
    if(ram_class_meta_field_type_21_is_repeated_MPORT_en & ram_class_meta_field_type_21_is_repeated_MPORT_mask) begin
      ram_class_meta_field_type_21_is_repeated[ram_class_meta_field_type_21_is_repeated_MPORT_addr] <=
        ram_class_meta_field_type_21_is_repeated_MPORT_data; // @[Decoupled.scala 218:16]
    end
    if(ram_class_meta_field_type_21_field_type_MPORT_en & ram_class_meta_field_type_21_field_type_MPORT_mask) begin
      ram_class_meta_field_type_21_field_type[ram_class_meta_field_type_21_field_type_MPORT_addr] <=
        ram_class_meta_field_type_21_field_type_MPORT_data; // @[Decoupled.scala 218:16]
    end
    if(ram_class_meta_field_type_21_sub_class_id_MPORT_en & ram_class_meta_field_type_21_sub_class_id_MPORT_mask) begin
      ram_class_meta_field_type_21_sub_class_id[ram_class_meta_field_type_21_sub_class_id_MPORT_addr] <=
        ram_class_meta_field_type_21_sub_class_id_MPORT_data; // @[Decoupled.scala 218:16]
    end
    if(ram_class_meta_field_type_22_is_repeated_MPORT_en & ram_class_meta_field_type_22_is_repeated_MPORT_mask) begin
      ram_class_meta_field_type_22_is_repeated[ram_class_meta_field_type_22_is_repeated_MPORT_addr] <=
        ram_class_meta_field_type_22_is_repeated_MPORT_data; // @[Decoupled.scala 218:16]
    end
    if(ram_class_meta_field_type_22_field_type_MPORT_en & ram_class_meta_field_type_22_field_type_MPORT_mask) begin
      ram_class_meta_field_type_22_field_type[ram_class_meta_field_type_22_field_type_MPORT_addr] <=
        ram_class_meta_field_type_22_field_type_MPORT_data; // @[Decoupled.scala 218:16]
    end
    if(ram_class_meta_field_type_22_sub_class_id_MPORT_en & ram_class_meta_field_type_22_sub_class_id_MPORT_mask) begin
      ram_class_meta_field_type_22_sub_class_id[ram_class_meta_field_type_22_sub_class_id_MPORT_addr] <=
        ram_class_meta_field_type_22_sub_class_id_MPORT_data; // @[Decoupled.scala 218:16]
    end
    if(ram_class_meta_field_type_23_is_repeated_MPORT_en & ram_class_meta_field_type_23_is_repeated_MPORT_mask) begin
      ram_class_meta_field_type_23_is_repeated[ram_class_meta_field_type_23_is_repeated_MPORT_addr] <=
        ram_class_meta_field_type_23_is_repeated_MPORT_data; // @[Decoupled.scala 218:16]
    end
    if(ram_class_meta_field_type_23_field_type_MPORT_en & ram_class_meta_field_type_23_field_type_MPORT_mask) begin
      ram_class_meta_field_type_23_field_type[ram_class_meta_field_type_23_field_type_MPORT_addr] <=
        ram_class_meta_field_type_23_field_type_MPORT_data; // @[Decoupled.scala 218:16]
    end
    if(ram_class_meta_field_type_23_sub_class_id_MPORT_en & ram_class_meta_field_type_23_sub_class_id_MPORT_mask) begin
      ram_class_meta_field_type_23_sub_class_id[ram_class_meta_field_type_23_sub_class_id_MPORT_addr] <=
        ram_class_meta_field_type_23_sub_class_id_MPORT_data; // @[Decoupled.scala 218:16]
    end
    if(ram_class_meta_field_type_24_is_repeated_MPORT_en & ram_class_meta_field_type_24_is_repeated_MPORT_mask) begin
      ram_class_meta_field_type_24_is_repeated[ram_class_meta_field_type_24_is_repeated_MPORT_addr] <=
        ram_class_meta_field_type_24_is_repeated_MPORT_data; // @[Decoupled.scala 218:16]
    end
    if(ram_class_meta_field_type_24_field_type_MPORT_en & ram_class_meta_field_type_24_field_type_MPORT_mask) begin
      ram_class_meta_field_type_24_field_type[ram_class_meta_field_type_24_field_type_MPORT_addr] <=
        ram_class_meta_field_type_24_field_type_MPORT_data; // @[Decoupled.scala 218:16]
    end
    if(ram_class_meta_field_type_24_sub_class_id_MPORT_en & ram_class_meta_field_type_24_sub_class_id_MPORT_mask) begin
      ram_class_meta_field_type_24_sub_class_id[ram_class_meta_field_type_24_sub_class_id_MPORT_addr] <=
        ram_class_meta_field_type_24_sub_class_id_MPORT_data; // @[Decoupled.scala 218:16]
    end
    if(ram_class_meta_field_type_25_is_repeated_MPORT_en & ram_class_meta_field_type_25_is_repeated_MPORT_mask) begin
      ram_class_meta_field_type_25_is_repeated[ram_class_meta_field_type_25_is_repeated_MPORT_addr] <=
        ram_class_meta_field_type_25_is_repeated_MPORT_data; // @[Decoupled.scala 218:16]
    end
    if(ram_class_meta_field_type_25_field_type_MPORT_en & ram_class_meta_field_type_25_field_type_MPORT_mask) begin
      ram_class_meta_field_type_25_field_type[ram_class_meta_field_type_25_field_type_MPORT_addr] <=
        ram_class_meta_field_type_25_field_type_MPORT_data; // @[Decoupled.scala 218:16]
    end
    if(ram_class_meta_field_type_25_sub_class_id_MPORT_en & ram_class_meta_field_type_25_sub_class_id_MPORT_mask) begin
      ram_class_meta_field_type_25_sub_class_id[ram_class_meta_field_type_25_sub_class_id_MPORT_addr] <=
        ram_class_meta_field_type_25_sub_class_id_MPORT_data; // @[Decoupled.scala 218:16]
    end
    if(ram_class_meta_field_type_26_is_repeated_MPORT_en & ram_class_meta_field_type_26_is_repeated_MPORT_mask) begin
      ram_class_meta_field_type_26_is_repeated[ram_class_meta_field_type_26_is_repeated_MPORT_addr] <=
        ram_class_meta_field_type_26_is_repeated_MPORT_data; // @[Decoupled.scala 218:16]
    end
    if(ram_class_meta_field_type_26_field_type_MPORT_en & ram_class_meta_field_type_26_field_type_MPORT_mask) begin
      ram_class_meta_field_type_26_field_type[ram_class_meta_field_type_26_field_type_MPORT_addr] <=
        ram_class_meta_field_type_26_field_type_MPORT_data; // @[Decoupled.scala 218:16]
    end
    if(ram_class_meta_field_type_26_sub_class_id_MPORT_en & ram_class_meta_field_type_26_sub_class_id_MPORT_mask) begin
      ram_class_meta_field_type_26_sub_class_id[ram_class_meta_field_type_26_sub_class_id_MPORT_addr] <=
        ram_class_meta_field_type_26_sub_class_id_MPORT_data; // @[Decoupled.scala 218:16]
    end
    if(ram_class_meta_field_type_27_is_repeated_MPORT_en & ram_class_meta_field_type_27_is_repeated_MPORT_mask) begin
      ram_class_meta_field_type_27_is_repeated[ram_class_meta_field_type_27_is_repeated_MPORT_addr] <=
        ram_class_meta_field_type_27_is_repeated_MPORT_data; // @[Decoupled.scala 218:16]
    end
    if(ram_class_meta_field_type_27_field_type_MPORT_en & ram_class_meta_field_type_27_field_type_MPORT_mask) begin
      ram_class_meta_field_type_27_field_type[ram_class_meta_field_type_27_field_type_MPORT_addr] <=
        ram_class_meta_field_type_27_field_type_MPORT_data; // @[Decoupled.scala 218:16]
    end
    if(ram_class_meta_field_type_27_sub_class_id_MPORT_en & ram_class_meta_field_type_27_sub_class_id_MPORT_mask) begin
      ram_class_meta_field_type_27_sub_class_id[ram_class_meta_field_type_27_sub_class_id_MPORT_addr] <=
        ram_class_meta_field_type_27_sub_class_id_MPORT_data; // @[Decoupled.scala 218:16]
    end
    if(ram_class_meta_field_type_28_is_repeated_MPORT_en & ram_class_meta_field_type_28_is_repeated_MPORT_mask) begin
      ram_class_meta_field_type_28_is_repeated[ram_class_meta_field_type_28_is_repeated_MPORT_addr] <=
        ram_class_meta_field_type_28_is_repeated_MPORT_data; // @[Decoupled.scala 218:16]
    end
    if(ram_class_meta_field_type_28_field_type_MPORT_en & ram_class_meta_field_type_28_field_type_MPORT_mask) begin
      ram_class_meta_field_type_28_field_type[ram_class_meta_field_type_28_field_type_MPORT_addr] <=
        ram_class_meta_field_type_28_field_type_MPORT_data; // @[Decoupled.scala 218:16]
    end
    if(ram_class_meta_field_type_28_sub_class_id_MPORT_en & ram_class_meta_field_type_28_sub_class_id_MPORT_mask) begin
      ram_class_meta_field_type_28_sub_class_id[ram_class_meta_field_type_28_sub_class_id_MPORT_addr] <=
        ram_class_meta_field_type_28_sub_class_id_MPORT_data; // @[Decoupled.scala 218:16]
    end
    if(ram_class_meta_field_type_29_is_repeated_MPORT_en & ram_class_meta_field_type_29_is_repeated_MPORT_mask) begin
      ram_class_meta_field_type_29_is_repeated[ram_class_meta_field_type_29_is_repeated_MPORT_addr] <=
        ram_class_meta_field_type_29_is_repeated_MPORT_data; // @[Decoupled.scala 218:16]
    end
    if(ram_class_meta_field_type_29_field_type_MPORT_en & ram_class_meta_field_type_29_field_type_MPORT_mask) begin
      ram_class_meta_field_type_29_field_type[ram_class_meta_field_type_29_field_type_MPORT_addr] <=
        ram_class_meta_field_type_29_field_type_MPORT_data; // @[Decoupled.scala 218:16]
    end
    if(ram_class_meta_field_type_29_sub_class_id_MPORT_en & ram_class_meta_field_type_29_sub_class_id_MPORT_mask) begin
      ram_class_meta_field_type_29_sub_class_id[ram_class_meta_field_type_29_sub_class_id_MPORT_addr] <=
        ram_class_meta_field_type_29_sub_class_id_MPORT_data; // @[Decoupled.scala 218:16]
    end
    if(ram_class_meta_field_type_30_is_repeated_MPORT_en & ram_class_meta_field_type_30_is_repeated_MPORT_mask) begin
      ram_class_meta_field_type_30_is_repeated[ram_class_meta_field_type_30_is_repeated_MPORT_addr] <=
        ram_class_meta_field_type_30_is_repeated_MPORT_data; // @[Decoupled.scala 218:16]
    end
    if(ram_class_meta_field_type_30_field_type_MPORT_en & ram_class_meta_field_type_30_field_type_MPORT_mask) begin
      ram_class_meta_field_type_30_field_type[ram_class_meta_field_type_30_field_type_MPORT_addr] <=
        ram_class_meta_field_type_30_field_type_MPORT_data; // @[Decoupled.scala 218:16]
    end
    if(ram_class_meta_field_type_30_sub_class_id_MPORT_en & ram_class_meta_field_type_30_sub_class_id_MPORT_mask) begin
      ram_class_meta_field_type_30_sub_class_id[ram_class_meta_field_type_30_sub_class_id_MPORT_addr] <=
        ram_class_meta_field_type_30_sub_class_id_MPORT_data; // @[Decoupled.scala 218:16]
    end
    if(ram_class_meta_field_type_31_is_repeated_MPORT_en & ram_class_meta_field_type_31_is_repeated_MPORT_mask) begin
      ram_class_meta_field_type_31_is_repeated[ram_class_meta_field_type_31_is_repeated_MPORT_addr] <=
        ram_class_meta_field_type_31_is_repeated_MPORT_data; // @[Decoupled.scala 218:16]
    end
    if(ram_class_meta_field_type_31_field_type_MPORT_en & ram_class_meta_field_type_31_field_type_MPORT_mask) begin
      ram_class_meta_field_type_31_field_type[ram_class_meta_field_type_31_field_type_MPORT_addr] <=
        ram_class_meta_field_type_31_field_type_MPORT_data; // @[Decoupled.scala 218:16]
    end
    if(ram_class_meta_field_type_31_sub_class_id_MPORT_en & ram_class_meta_field_type_31_sub_class_id_MPORT_mask) begin
      ram_class_meta_field_type_31_sub_class_id[ram_class_meta_field_type_31_sub_class_id_MPORT_addr] <=
        ram_class_meta_field_type_31_sub_class_id_MPORT_data; // @[Decoupled.scala 218:16]
    end
    if(ram_class_meta_field_type_32_is_repeated_MPORT_en & ram_class_meta_field_type_32_is_repeated_MPORT_mask) begin
      ram_class_meta_field_type_32_is_repeated[ram_class_meta_field_type_32_is_repeated_MPORT_addr] <=
        ram_class_meta_field_type_32_is_repeated_MPORT_data; // @[Decoupled.scala 218:16]
    end
    if(ram_class_meta_field_type_32_field_type_MPORT_en & ram_class_meta_field_type_32_field_type_MPORT_mask) begin
      ram_class_meta_field_type_32_field_type[ram_class_meta_field_type_32_field_type_MPORT_addr] <=
        ram_class_meta_field_type_32_field_type_MPORT_data; // @[Decoupled.scala 218:16]
    end
    if(ram_class_meta_field_type_32_sub_class_id_MPORT_en & ram_class_meta_field_type_32_sub_class_id_MPORT_mask) begin
      ram_class_meta_field_type_32_sub_class_id[ram_class_meta_field_type_32_sub_class_id_MPORT_addr] <=
        ram_class_meta_field_type_32_sub_class_id_MPORT_data; // @[Decoupled.scala 218:16]
    end
    if (reset) begin // @[Counter.scala 60:40]
      enq_ptr_value <= 3'h0; // @[Counter.scala 60:40]
    end else if (do_enq) begin // @[Decoupled.scala 229:17]
      enq_ptr_value <= _value_T_1; // @[Counter.scala 76:15]
    end
    if (reset) begin // @[Counter.scala 60:40]
      deq_ptr_value <= 3'h0; // @[Counter.scala 60:40]
    end else if (do_deq) begin // @[Decoupled.scala 233:17]
      deq_ptr_value <= _value_T_3; // @[Counter.scala 76:15]
    end
    if (reset) begin // @[Decoupled.scala 221:27]
      maybe_full <= 1'h0; // @[Decoupled.scala 221:27]
    end else if (do_enq != do_deq) begin // @[Decoupled.scala 236:28]
      maybe_full <= do_enq; // @[Decoupled.scala 237:16]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 8; initvar = initvar+1)
    ram_class_meta_max_field_num[initvar] = _RAND_0[7:0];
  _RAND_1 = {1{`RANDOM}};
  for (initvar = 0; initvar < 8; initvar = initvar+1)
    ram_class_meta_field_type_0_is_repeated[initvar] = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  for (initvar = 0; initvar < 8; initvar = initvar+1)
    ram_class_meta_field_type_0_field_type[initvar] = _RAND_2[4:0];
  _RAND_3 = {1{`RANDOM}};
  for (initvar = 0; initvar < 8; initvar = initvar+1)
    ram_class_meta_field_type_0_sub_class_id[initvar] = _RAND_3[15:0];
  _RAND_4 = {1{`RANDOM}};
  for (initvar = 0; initvar < 8; initvar = initvar+1)
    ram_class_meta_field_type_1_is_repeated[initvar] = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  for (initvar = 0; initvar < 8; initvar = initvar+1)
    ram_class_meta_field_type_1_field_type[initvar] = _RAND_5[4:0];
  _RAND_6 = {1{`RANDOM}};
  for (initvar = 0; initvar < 8; initvar = initvar+1)
    ram_class_meta_field_type_1_sub_class_id[initvar] = _RAND_6[15:0];
  _RAND_7 = {1{`RANDOM}};
  for (initvar = 0; initvar < 8; initvar = initvar+1)
    ram_class_meta_field_type_2_is_repeated[initvar] = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  for (initvar = 0; initvar < 8; initvar = initvar+1)
    ram_class_meta_field_type_2_field_type[initvar] = _RAND_8[4:0];
  _RAND_9 = {1{`RANDOM}};
  for (initvar = 0; initvar < 8; initvar = initvar+1)
    ram_class_meta_field_type_2_sub_class_id[initvar] = _RAND_9[15:0];
  _RAND_10 = {1{`RANDOM}};
  for (initvar = 0; initvar < 8; initvar = initvar+1)
    ram_class_meta_field_type_3_is_repeated[initvar] = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  for (initvar = 0; initvar < 8; initvar = initvar+1)
    ram_class_meta_field_type_3_field_type[initvar] = _RAND_11[4:0];
  _RAND_12 = {1{`RANDOM}};
  for (initvar = 0; initvar < 8; initvar = initvar+1)
    ram_class_meta_field_type_3_sub_class_id[initvar] = _RAND_12[15:0];
  _RAND_13 = {1{`RANDOM}};
  for (initvar = 0; initvar < 8; initvar = initvar+1)
    ram_class_meta_field_type_4_is_repeated[initvar] = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  for (initvar = 0; initvar < 8; initvar = initvar+1)
    ram_class_meta_field_type_4_field_type[initvar] = _RAND_14[4:0];
  _RAND_15 = {1{`RANDOM}};
  for (initvar = 0; initvar < 8; initvar = initvar+1)
    ram_class_meta_field_type_4_sub_class_id[initvar] = _RAND_15[15:0];
  _RAND_16 = {1{`RANDOM}};
  for (initvar = 0; initvar < 8; initvar = initvar+1)
    ram_class_meta_field_type_5_is_repeated[initvar] = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  for (initvar = 0; initvar < 8; initvar = initvar+1)
    ram_class_meta_field_type_5_field_type[initvar] = _RAND_17[4:0];
  _RAND_18 = {1{`RANDOM}};
  for (initvar = 0; initvar < 8; initvar = initvar+1)
    ram_class_meta_field_type_5_sub_class_id[initvar] = _RAND_18[15:0];
  _RAND_19 = {1{`RANDOM}};
  for (initvar = 0; initvar < 8; initvar = initvar+1)
    ram_class_meta_field_type_6_is_repeated[initvar] = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  for (initvar = 0; initvar < 8; initvar = initvar+1)
    ram_class_meta_field_type_6_field_type[initvar] = _RAND_20[4:0];
  _RAND_21 = {1{`RANDOM}};
  for (initvar = 0; initvar < 8; initvar = initvar+1)
    ram_class_meta_field_type_6_sub_class_id[initvar] = _RAND_21[15:0];
  _RAND_22 = {1{`RANDOM}};
  for (initvar = 0; initvar < 8; initvar = initvar+1)
    ram_class_meta_field_type_7_is_repeated[initvar] = _RAND_22[0:0];
  _RAND_23 = {1{`RANDOM}};
  for (initvar = 0; initvar < 8; initvar = initvar+1)
    ram_class_meta_field_type_7_field_type[initvar] = _RAND_23[4:0];
  _RAND_24 = {1{`RANDOM}};
  for (initvar = 0; initvar < 8; initvar = initvar+1)
    ram_class_meta_field_type_7_sub_class_id[initvar] = _RAND_24[15:0];
  _RAND_25 = {1{`RANDOM}};
  for (initvar = 0; initvar < 8; initvar = initvar+1)
    ram_class_meta_field_type_8_is_repeated[initvar] = _RAND_25[0:0];
  _RAND_26 = {1{`RANDOM}};
  for (initvar = 0; initvar < 8; initvar = initvar+1)
    ram_class_meta_field_type_8_field_type[initvar] = _RAND_26[4:0];
  _RAND_27 = {1{`RANDOM}};
  for (initvar = 0; initvar < 8; initvar = initvar+1)
    ram_class_meta_field_type_8_sub_class_id[initvar] = _RAND_27[15:0];
  _RAND_28 = {1{`RANDOM}};
  for (initvar = 0; initvar < 8; initvar = initvar+1)
    ram_class_meta_field_type_9_is_repeated[initvar] = _RAND_28[0:0];
  _RAND_29 = {1{`RANDOM}};
  for (initvar = 0; initvar < 8; initvar = initvar+1)
    ram_class_meta_field_type_9_field_type[initvar] = _RAND_29[4:0];
  _RAND_30 = {1{`RANDOM}};
  for (initvar = 0; initvar < 8; initvar = initvar+1)
    ram_class_meta_field_type_9_sub_class_id[initvar] = _RAND_30[15:0];
  _RAND_31 = {1{`RANDOM}};
  for (initvar = 0; initvar < 8; initvar = initvar+1)
    ram_class_meta_field_type_10_is_repeated[initvar] = _RAND_31[0:0];
  _RAND_32 = {1{`RANDOM}};
  for (initvar = 0; initvar < 8; initvar = initvar+1)
    ram_class_meta_field_type_10_field_type[initvar] = _RAND_32[4:0];
  _RAND_33 = {1{`RANDOM}};
  for (initvar = 0; initvar < 8; initvar = initvar+1)
    ram_class_meta_field_type_10_sub_class_id[initvar] = _RAND_33[15:0];
  _RAND_34 = {1{`RANDOM}};
  for (initvar = 0; initvar < 8; initvar = initvar+1)
    ram_class_meta_field_type_11_is_repeated[initvar] = _RAND_34[0:0];
  _RAND_35 = {1{`RANDOM}};
  for (initvar = 0; initvar < 8; initvar = initvar+1)
    ram_class_meta_field_type_11_field_type[initvar] = _RAND_35[4:0];
  _RAND_36 = {1{`RANDOM}};
  for (initvar = 0; initvar < 8; initvar = initvar+1)
    ram_class_meta_field_type_11_sub_class_id[initvar] = _RAND_36[15:0];
  _RAND_37 = {1{`RANDOM}};
  for (initvar = 0; initvar < 8; initvar = initvar+1)
    ram_class_meta_field_type_12_is_repeated[initvar] = _RAND_37[0:0];
  _RAND_38 = {1{`RANDOM}};
  for (initvar = 0; initvar < 8; initvar = initvar+1)
    ram_class_meta_field_type_12_field_type[initvar] = _RAND_38[4:0];
  _RAND_39 = {1{`RANDOM}};
  for (initvar = 0; initvar < 8; initvar = initvar+1)
    ram_class_meta_field_type_12_sub_class_id[initvar] = _RAND_39[15:0];
  _RAND_40 = {1{`RANDOM}};
  for (initvar = 0; initvar < 8; initvar = initvar+1)
    ram_class_meta_field_type_13_is_repeated[initvar] = _RAND_40[0:0];
  _RAND_41 = {1{`RANDOM}};
  for (initvar = 0; initvar < 8; initvar = initvar+1)
    ram_class_meta_field_type_13_field_type[initvar] = _RAND_41[4:0];
  _RAND_42 = {1{`RANDOM}};
  for (initvar = 0; initvar < 8; initvar = initvar+1)
    ram_class_meta_field_type_13_sub_class_id[initvar] = _RAND_42[15:0];
  _RAND_43 = {1{`RANDOM}};
  for (initvar = 0; initvar < 8; initvar = initvar+1)
    ram_class_meta_field_type_14_is_repeated[initvar] = _RAND_43[0:0];
  _RAND_44 = {1{`RANDOM}};
  for (initvar = 0; initvar < 8; initvar = initvar+1)
    ram_class_meta_field_type_14_field_type[initvar] = _RAND_44[4:0];
  _RAND_45 = {1{`RANDOM}};
  for (initvar = 0; initvar < 8; initvar = initvar+1)
    ram_class_meta_field_type_14_sub_class_id[initvar] = _RAND_45[15:0];
  _RAND_46 = {1{`RANDOM}};
  for (initvar = 0; initvar < 8; initvar = initvar+1)
    ram_class_meta_field_type_15_is_repeated[initvar] = _RAND_46[0:0];
  _RAND_47 = {1{`RANDOM}};
  for (initvar = 0; initvar < 8; initvar = initvar+1)
    ram_class_meta_field_type_15_field_type[initvar] = _RAND_47[4:0];
  _RAND_48 = {1{`RANDOM}};
  for (initvar = 0; initvar < 8; initvar = initvar+1)
    ram_class_meta_field_type_15_sub_class_id[initvar] = _RAND_48[15:0];
  _RAND_49 = {1{`RANDOM}};
  for (initvar = 0; initvar < 8; initvar = initvar+1)
    ram_class_meta_field_type_16_is_repeated[initvar] = _RAND_49[0:0];
  _RAND_50 = {1{`RANDOM}};
  for (initvar = 0; initvar < 8; initvar = initvar+1)
    ram_class_meta_field_type_16_field_type[initvar] = _RAND_50[4:0];
  _RAND_51 = {1{`RANDOM}};
  for (initvar = 0; initvar < 8; initvar = initvar+1)
    ram_class_meta_field_type_16_sub_class_id[initvar] = _RAND_51[15:0];
  _RAND_52 = {1{`RANDOM}};
  for (initvar = 0; initvar < 8; initvar = initvar+1)
    ram_class_meta_field_type_17_is_repeated[initvar] = _RAND_52[0:0];
  _RAND_53 = {1{`RANDOM}};
  for (initvar = 0; initvar < 8; initvar = initvar+1)
    ram_class_meta_field_type_17_field_type[initvar] = _RAND_53[4:0];
  _RAND_54 = {1{`RANDOM}};
  for (initvar = 0; initvar < 8; initvar = initvar+1)
    ram_class_meta_field_type_17_sub_class_id[initvar] = _RAND_54[15:0];
  _RAND_55 = {1{`RANDOM}};
  for (initvar = 0; initvar < 8; initvar = initvar+1)
    ram_class_meta_field_type_18_is_repeated[initvar] = _RAND_55[0:0];
  _RAND_56 = {1{`RANDOM}};
  for (initvar = 0; initvar < 8; initvar = initvar+1)
    ram_class_meta_field_type_18_field_type[initvar] = _RAND_56[4:0];
  _RAND_57 = {1{`RANDOM}};
  for (initvar = 0; initvar < 8; initvar = initvar+1)
    ram_class_meta_field_type_18_sub_class_id[initvar] = _RAND_57[15:0];
  _RAND_58 = {1{`RANDOM}};
  for (initvar = 0; initvar < 8; initvar = initvar+1)
    ram_class_meta_field_type_19_is_repeated[initvar] = _RAND_58[0:0];
  _RAND_59 = {1{`RANDOM}};
  for (initvar = 0; initvar < 8; initvar = initvar+1)
    ram_class_meta_field_type_19_field_type[initvar] = _RAND_59[4:0];
  _RAND_60 = {1{`RANDOM}};
  for (initvar = 0; initvar < 8; initvar = initvar+1)
    ram_class_meta_field_type_19_sub_class_id[initvar] = _RAND_60[15:0];
  _RAND_61 = {1{`RANDOM}};
  for (initvar = 0; initvar < 8; initvar = initvar+1)
    ram_class_meta_field_type_20_is_repeated[initvar] = _RAND_61[0:0];
  _RAND_62 = {1{`RANDOM}};
  for (initvar = 0; initvar < 8; initvar = initvar+1)
    ram_class_meta_field_type_20_field_type[initvar] = _RAND_62[4:0];
  _RAND_63 = {1{`RANDOM}};
  for (initvar = 0; initvar < 8; initvar = initvar+1)
    ram_class_meta_field_type_20_sub_class_id[initvar] = _RAND_63[15:0];
  _RAND_64 = {1{`RANDOM}};
  for (initvar = 0; initvar < 8; initvar = initvar+1)
    ram_class_meta_field_type_21_is_repeated[initvar] = _RAND_64[0:0];
  _RAND_65 = {1{`RANDOM}};
  for (initvar = 0; initvar < 8; initvar = initvar+1)
    ram_class_meta_field_type_21_field_type[initvar] = _RAND_65[4:0];
  _RAND_66 = {1{`RANDOM}};
  for (initvar = 0; initvar < 8; initvar = initvar+1)
    ram_class_meta_field_type_21_sub_class_id[initvar] = _RAND_66[15:0];
  _RAND_67 = {1{`RANDOM}};
  for (initvar = 0; initvar < 8; initvar = initvar+1)
    ram_class_meta_field_type_22_is_repeated[initvar] = _RAND_67[0:0];
  _RAND_68 = {1{`RANDOM}};
  for (initvar = 0; initvar < 8; initvar = initvar+1)
    ram_class_meta_field_type_22_field_type[initvar] = _RAND_68[4:0];
  _RAND_69 = {1{`RANDOM}};
  for (initvar = 0; initvar < 8; initvar = initvar+1)
    ram_class_meta_field_type_22_sub_class_id[initvar] = _RAND_69[15:0];
  _RAND_70 = {1{`RANDOM}};
  for (initvar = 0; initvar < 8; initvar = initvar+1)
    ram_class_meta_field_type_23_is_repeated[initvar] = _RAND_70[0:0];
  _RAND_71 = {1{`RANDOM}};
  for (initvar = 0; initvar < 8; initvar = initvar+1)
    ram_class_meta_field_type_23_field_type[initvar] = _RAND_71[4:0];
  _RAND_72 = {1{`RANDOM}};
  for (initvar = 0; initvar < 8; initvar = initvar+1)
    ram_class_meta_field_type_23_sub_class_id[initvar] = _RAND_72[15:0];
  _RAND_73 = {1{`RANDOM}};
  for (initvar = 0; initvar < 8; initvar = initvar+1)
    ram_class_meta_field_type_24_is_repeated[initvar] = _RAND_73[0:0];
  _RAND_74 = {1{`RANDOM}};
  for (initvar = 0; initvar < 8; initvar = initvar+1)
    ram_class_meta_field_type_24_field_type[initvar] = _RAND_74[4:0];
  _RAND_75 = {1{`RANDOM}};
  for (initvar = 0; initvar < 8; initvar = initvar+1)
    ram_class_meta_field_type_24_sub_class_id[initvar] = _RAND_75[15:0];
  _RAND_76 = {1{`RANDOM}};
  for (initvar = 0; initvar < 8; initvar = initvar+1)
    ram_class_meta_field_type_25_is_repeated[initvar] = _RAND_76[0:0];
  _RAND_77 = {1{`RANDOM}};
  for (initvar = 0; initvar < 8; initvar = initvar+1)
    ram_class_meta_field_type_25_field_type[initvar] = _RAND_77[4:0];
  _RAND_78 = {1{`RANDOM}};
  for (initvar = 0; initvar < 8; initvar = initvar+1)
    ram_class_meta_field_type_25_sub_class_id[initvar] = _RAND_78[15:0];
  _RAND_79 = {1{`RANDOM}};
  for (initvar = 0; initvar < 8; initvar = initvar+1)
    ram_class_meta_field_type_26_is_repeated[initvar] = _RAND_79[0:0];
  _RAND_80 = {1{`RANDOM}};
  for (initvar = 0; initvar < 8; initvar = initvar+1)
    ram_class_meta_field_type_26_field_type[initvar] = _RAND_80[4:0];
  _RAND_81 = {1{`RANDOM}};
  for (initvar = 0; initvar < 8; initvar = initvar+1)
    ram_class_meta_field_type_26_sub_class_id[initvar] = _RAND_81[15:0];
  _RAND_82 = {1{`RANDOM}};
  for (initvar = 0; initvar < 8; initvar = initvar+1)
    ram_class_meta_field_type_27_is_repeated[initvar] = _RAND_82[0:0];
  _RAND_83 = {1{`RANDOM}};
  for (initvar = 0; initvar < 8; initvar = initvar+1)
    ram_class_meta_field_type_27_field_type[initvar] = _RAND_83[4:0];
  _RAND_84 = {1{`RANDOM}};
  for (initvar = 0; initvar < 8; initvar = initvar+1)
    ram_class_meta_field_type_27_sub_class_id[initvar] = _RAND_84[15:0];
  _RAND_85 = {1{`RANDOM}};
  for (initvar = 0; initvar < 8; initvar = initvar+1)
    ram_class_meta_field_type_28_is_repeated[initvar] = _RAND_85[0:0];
  _RAND_86 = {1{`RANDOM}};
  for (initvar = 0; initvar < 8; initvar = initvar+1)
    ram_class_meta_field_type_28_field_type[initvar] = _RAND_86[4:0];
  _RAND_87 = {1{`RANDOM}};
  for (initvar = 0; initvar < 8; initvar = initvar+1)
    ram_class_meta_field_type_28_sub_class_id[initvar] = _RAND_87[15:0];
  _RAND_88 = {1{`RANDOM}};
  for (initvar = 0; initvar < 8; initvar = initvar+1)
    ram_class_meta_field_type_29_is_repeated[initvar] = _RAND_88[0:0];
  _RAND_89 = {1{`RANDOM}};
  for (initvar = 0; initvar < 8; initvar = initvar+1)
    ram_class_meta_field_type_29_field_type[initvar] = _RAND_89[4:0];
  _RAND_90 = {1{`RANDOM}};
  for (initvar = 0; initvar < 8; initvar = initvar+1)
    ram_class_meta_field_type_29_sub_class_id[initvar] = _RAND_90[15:0];
  _RAND_91 = {1{`RANDOM}};
  for (initvar = 0; initvar < 8; initvar = initvar+1)
    ram_class_meta_field_type_30_is_repeated[initvar] = _RAND_91[0:0];
  _RAND_92 = {1{`RANDOM}};
  for (initvar = 0; initvar < 8; initvar = initvar+1)
    ram_class_meta_field_type_30_field_type[initvar] = _RAND_92[4:0];
  _RAND_93 = {1{`RANDOM}};
  for (initvar = 0; initvar < 8; initvar = initvar+1)
    ram_class_meta_field_type_30_sub_class_id[initvar] = _RAND_93[15:0];
  _RAND_94 = {1{`RANDOM}};
  for (initvar = 0; initvar < 8; initvar = initvar+1)
    ram_class_meta_field_type_31_is_repeated[initvar] = _RAND_94[0:0];
  _RAND_95 = {1{`RANDOM}};
  for (initvar = 0; initvar < 8; initvar = initvar+1)
    ram_class_meta_field_type_31_field_type[initvar] = _RAND_95[4:0];
  _RAND_96 = {1{`RANDOM}};
  for (initvar = 0; initvar < 8; initvar = initvar+1)
    ram_class_meta_field_type_31_sub_class_id[initvar] = _RAND_96[15:0];
  _RAND_97 = {1{`RANDOM}};
  for (initvar = 0; initvar < 8; initvar = initvar+1)
    ram_class_meta_field_type_32_is_repeated[initvar] = _RAND_97[0:0];
  _RAND_98 = {1{`RANDOM}};
  for (initvar = 0; initvar < 8; initvar = initvar+1)
    ram_class_meta_field_type_32_field_type[initvar] = _RAND_98[4:0];
  _RAND_99 = {1{`RANDOM}};
  for (initvar = 0; initvar < 8; initvar = initvar+1)
    ram_class_meta_field_type_32_sub_class_id[initvar] = _RAND_99[15:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_100 = {1{`RANDOM}};
  enq_ptr_value = _RAND_100[2:0];
  _RAND_101 = {1{`RANDOM}};
  deq_ptr_value = _RAND_101[2:0];
  _RAND_102 = {1{`RANDOM}};
  maybe_full = _RAND_102[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module XQueue_3(
  input         clock,
  input         reset,
  input         io_in_valid,
  input  [7:0]  io_in_bits_class_meta_max_field_num,
  input         io_in_bits_class_meta_field_type_0_is_repeated,
  input  [4:0]  io_in_bits_class_meta_field_type_0_field_type,
  input  [15:0] io_in_bits_class_meta_field_type_0_sub_class_id,
  input         io_in_bits_class_meta_field_type_1_is_repeated,
  input  [4:0]  io_in_bits_class_meta_field_type_1_field_type,
  input  [15:0] io_in_bits_class_meta_field_type_1_sub_class_id,
  input         io_in_bits_class_meta_field_type_2_is_repeated,
  input  [4:0]  io_in_bits_class_meta_field_type_2_field_type,
  input  [15:0] io_in_bits_class_meta_field_type_2_sub_class_id,
  input         io_in_bits_class_meta_field_type_3_is_repeated,
  input  [4:0]  io_in_bits_class_meta_field_type_3_field_type,
  input  [15:0] io_in_bits_class_meta_field_type_3_sub_class_id,
  input         io_in_bits_class_meta_field_type_4_is_repeated,
  input  [4:0]  io_in_bits_class_meta_field_type_4_field_type,
  input  [15:0] io_in_bits_class_meta_field_type_4_sub_class_id,
  input         io_in_bits_class_meta_field_type_5_is_repeated,
  input  [4:0]  io_in_bits_class_meta_field_type_5_field_type,
  input  [15:0] io_in_bits_class_meta_field_type_5_sub_class_id,
  input         io_in_bits_class_meta_field_type_6_is_repeated,
  input  [4:0]  io_in_bits_class_meta_field_type_6_field_type,
  input  [15:0] io_in_bits_class_meta_field_type_6_sub_class_id,
  input         io_in_bits_class_meta_field_type_7_is_repeated,
  input  [4:0]  io_in_bits_class_meta_field_type_7_field_type,
  input  [15:0] io_in_bits_class_meta_field_type_7_sub_class_id,
  input         io_in_bits_class_meta_field_type_8_is_repeated,
  input  [4:0]  io_in_bits_class_meta_field_type_8_field_type,
  input  [15:0] io_in_bits_class_meta_field_type_8_sub_class_id,
  input         io_in_bits_class_meta_field_type_9_is_repeated,
  input  [4:0]  io_in_bits_class_meta_field_type_9_field_type,
  input  [15:0] io_in_bits_class_meta_field_type_9_sub_class_id,
  input         io_in_bits_class_meta_field_type_10_is_repeated,
  input  [4:0]  io_in_bits_class_meta_field_type_10_field_type,
  input  [15:0] io_in_bits_class_meta_field_type_10_sub_class_id,
  input         io_in_bits_class_meta_field_type_11_is_repeated,
  input  [4:0]  io_in_bits_class_meta_field_type_11_field_type,
  input  [15:0] io_in_bits_class_meta_field_type_11_sub_class_id,
  input         io_in_bits_class_meta_field_type_12_is_repeated,
  input  [4:0]  io_in_bits_class_meta_field_type_12_field_type,
  input  [15:0] io_in_bits_class_meta_field_type_12_sub_class_id,
  input         io_in_bits_class_meta_field_type_13_is_repeated,
  input  [4:0]  io_in_bits_class_meta_field_type_13_field_type,
  input  [15:0] io_in_bits_class_meta_field_type_13_sub_class_id,
  input         io_in_bits_class_meta_field_type_14_is_repeated,
  input  [4:0]  io_in_bits_class_meta_field_type_14_field_type,
  input  [15:0] io_in_bits_class_meta_field_type_14_sub_class_id,
  input         io_in_bits_class_meta_field_type_15_is_repeated,
  input  [4:0]  io_in_bits_class_meta_field_type_15_field_type,
  input  [15:0] io_in_bits_class_meta_field_type_15_sub_class_id,
  input         io_in_bits_class_meta_field_type_16_is_repeated,
  input  [4:0]  io_in_bits_class_meta_field_type_16_field_type,
  input  [15:0] io_in_bits_class_meta_field_type_16_sub_class_id,
  input         io_in_bits_class_meta_field_type_17_is_repeated,
  input  [4:0]  io_in_bits_class_meta_field_type_17_field_type,
  input  [15:0] io_in_bits_class_meta_field_type_17_sub_class_id,
  input         io_in_bits_class_meta_field_type_18_is_repeated,
  input  [4:0]  io_in_bits_class_meta_field_type_18_field_type,
  input  [15:0] io_in_bits_class_meta_field_type_18_sub_class_id,
  input         io_in_bits_class_meta_field_type_19_is_repeated,
  input  [4:0]  io_in_bits_class_meta_field_type_19_field_type,
  input  [15:0] io_in_bits_class_meta_field_type_19_sub_class_id,
  input         io_in_bits_class_meta_field_type_20_is_repeated,
  input  [4:0]  io_in_bits_class_meta_field_type_20_field_type,
  input  [15:0] io_in_bits_class_meta_field_type_20_sub_class_id,
  input         io_in_bits_class_meta_field_type_21_is_repeated,
  input  [4:0]  io_in_bits_class_meta_field_type_21_field_type,
  input  [15:0] io_in_bits_class_meta_field_type_21_sub_class_id,
  input         io_in_bits_class_meta_field_type_22_is_repeated,
  input  [4:0]  io_in_bits_class_meta_field_type_22_field_type,
  input  [15:0] io_in_bits_class_meta_field_type_22_sub_class_id,
  input         io_in_bits_class_meta_field_type_23_is_repeated,
  input  [4:0]  io_in_bits_class_meta_field_type_23_field_type,
  input  [15:0] io_in_bits_class_meta_field_type_23_sub_class_id,
  input         io_in_bits_class_meta_field_type_24_is_repeated,
  input  [4:0]  io_in_bits_class_meta_field_type_24_field_type,
  input  [15:0] io_in_bits_class_meta_field_type_24_sub_class_id,
  input         io_in_bits_class_meta_field_type_25_is_repeated,
  input  [4:0]  io_in_bits_class_meta_field_type_25_field_type,
  input  [15:0] io_in_bits_class_meta_field_type_25_sub_class_id,
  input         io_in_bits_class_meta_field_type_26_is_repeated,
  input  [4:0]  io_in_bits_class_meta_field_type_26_field_type,
  input  [15:0] io_in_bits_class_meta_field_type_26_sub_class_id,
  input         io_in_bits_class_meta_field_type_27_is_repeated,
  input  [4:0]  io_in_bits_class_meta_field_type_27_field_type,
  input  [15:0] io_in_bits_class_meta_field_type_27_sub_class_id,
  input         io_in_bits_class_meta_field_type_28_is_repeated,
  input  [4:0]  io_in_bits_class_meta_field_type_28_field_type,
  input  [15:0] io_in_bits_class_meta_field_type_28_sub_class_id,
  input         io_in_bits_class_meta_field_type_29_is_repeated,
  input  [4:0]  io_in_bits_class_meta_field_type_29_field_type,
  input  [15:0] io_in_bits_class_meta_field_type_29_sub_class_id,
  input         io_in_bits_class_meta_field_type_30_is_repeated,
  input  [4:0]  io_in_bits_class_meta_field_type_30_field_type,
  input  [15:0] io_in_bits_class_meta_field_type_30_sub_class_id,
  input         io_in_bits_class_meta_field_type_31_is_repeated,
  input  [4:0]  io_in_bits_class_meta_field_type_31_field_type,
  input  [15:0] io_in_bits_class_meta_field_type_31_sub_class_id,
  input         io_in_bits_class_meta_field_type_32_is_repeated,
  input  [4:0]  io_in_bits_class_meta_field_type_32_field_type,
  input  [15:0] io_in_bits_class_meta_field_type_32_sub_class_id,
  input         io_out_ready,
  output        io_out_valid,
  output [7:0]  io_out_bits_class_meta_max_field_num,
  output        io_out_bits_class_meta_field_type_0_is_repeated,
  output [4:0]  io_out_bits_class_meta_field_type_0_field_type,
  output [15:0] io_out_bits_class_meta_field_type_0_sub_class_id,
  output        io_out_bits_class_meta_field_type_1_is_repeated,
  output [4:0]  io_out_bits_class_meta_field_type_1_field_type,
  output [15:0] io_out_bits_class_meta_field_type_1_sub_class_id,
  output        io_out_bits_class_meta_field_type_2_is_repeated,
  output [4:0]  io_out_bits_class_meta_field_type_2_field_type,
  output [15:0] io_out_bits_class_meta_field_type_2_sub_class_id,
  output        io_out_bits_class_meta_field_type_3_is_repeated,
  output [4:0]  io_out_bits_class_meta_field_type_3_field_type,
  output [15:0] io_out_bits_class_meta_field_type_3_sub_class_id,
  output        io_out_bits_class_meta_field_type_4_is_repeated,
  output [4:0]  io_out_bits_class_meta_field_type_4_field_type,
  output [15:0] io_out_bits_class_meta_field_type_4_sub_class_id,
  output        io_out_bits_class_meta_field_type_5_is_repeated,
  output [4:0]  io_out_bits_class_meta_field_type_5_field_type,
  output [15:0] io_out_bits_class_meta_field_type_5_sub_class_id,
  output        io_out_bits_class_meta_field_type_6_is_repeated,
  output [4:0]  io_out_bits_class_meta_field_type_6_field_type,
  output [15:0] io_out_bits_class_meta_field_type_6_sub_class_id,
  output        io_out_bits_class_meta_field_type_7_is_repeated,
  output [4:0]  io_out_bits_class_meta_field_type_7_field_type,
  output [15:0] io_out_bits_class_meta_field_type_7_sub_class_id,
  output        io_out_bits_class_meta_field_type_8_is_repeated,
  output [4:0]  io_out_bits_class_meta_field_type_8_field_type,
  output [15:0] io_out_bits_class_meta_field_type_8_sub_class_id,
  output        io_out_bits_class_meta_field_type_9_is_repeated,
  output [4:0]  io_out_bits_class_meta_field_type_9_field_type,
  output [15:0] io_out_bits_class_meta_field_type_9_sub_class_id,
  output        io_out_bits_class_meta_field_type_10_is_repeated,
  output [4:0]  io_out_bits_class_meta_field_type_10_field_type,
  output [15:0] io_out_bits_class_meta_field_type_10_sub_class_id,
  output        io_out_bits_class_meta_field_type_11_is_repeated,
  output [4:0]  io_out_bits_class_meta_field_type_11_field_type,
  output [15:0] io_out_bits_class_meta_field_type_11_sub_class_id,
  output        io_out_bits_class_meta_field_type_12_is_repeated,
  output [4:0]  io_out_bits_class_meta_field_type_12_field_type,
  output [15:0] io_out_bits_class_meta_field_type_12_sub_class_id,
  output        io_out_bits_class_meta_field_type_13_is_repeated,
  output [4:0]  io_out_bits_class_meta_field_type_13_field_type,
  output [15:0] io_out_bits_class_meta_field_type_13_sub_class_id,
  output        io_out_bits_class_meta_field_type_14_is_repeated,
  output [4:0]  io_out_bits_class_meta_field_type_14_field_type,
  output [15:0] io_out_bits_class_meta_field_type_14_sub_class_id,
  output        io_out_bits_class_meta_field_type_15_is_repeated,
  output [4:0]  io_out_bits_class_meta_field_type_15_field_type,
  output [15:0] io_out_bits_class_meta_field_type_15_sub_class_id,
  output        io_out_bits_class_meta_field_type_16_is_repeated,
  output [4:0]  io_out_bits_class_meta_field_type_16_field_type,
  output [15:0] io_out_bits_class_meta_field_type_16_sub_class_id,
  output        io_out_bits_class_meta_field_type_17_is_repeated,
  output [4:0]  io_out_bits_class_meta_field_type_17_field_type,
  output [15:0] io_out_bits_class_meta_field_type_17_sub_class_id,
  output        io_out_bits_class_meta_field_type_18_is_repeated,
  output [4:0]  io_out_bits_class_meta_field_type_18_field_type,
  output [15:0] io_out_bits_class_meta_field_type_18_sub_class_id,
  output        io_out_bits_class_meta_field_type_19_is_repeated,
  output [4:0]  io_out_bits_class_meta_field_type_19_field_type,
  output [15:0] io_out_bits_class_meta_field_type_19_sub_class_id,
  output        io_out_bits_class_meta_field_type_20_is_repeated,
  output [4:0]  io_out_bits_class_meta_field_type_20_field_type,
  output [15:0] io_out_bits_class_meta_field_type_20_sub_class_id,
  output        io_out_bits_class_meta_field_type_21_is_repeated,
  output [4:0]  io_out_bits_class_meta_field_type_21_field_type,
  output [15:0] io_out_bits_class_meta_field_type_21_sub_class_id,
  output        io_out_bits_class_meta_field_type_22_is_repeated,
  output [4:0]  io_out_bits_class_meta_field_type_22_field_type,
  output [15:0] io_out_bits_class_meta_field_type_22_sub_class_id,
  output        io_out_bits_class_meta_field_type_23_is_repeated,
  output [4:0]  io_out_bits_class_meta_field_type_23_field_type,
  output [15:0] io_out_bits_class_meta_field_type_23_sub_class_id,
  output        io_out_bits_class_meta_field_type_24_is_repeated,
  output [4:0]  io_out_bits_class_meta_field_type_24_field_type,
  output [15:0] io_out_bits_class_meta_field_type_24_sub_class_id,
  output        io_out_bits_class_meta_field_type_25_is_repeated,
  output [4:0]  io_out_bits_class_meta_field_type_25_field_type,
  output [15:0] io_out_bits_class_meta_field_type_25_sub_class_id,
  output        io_out_bits_class_meta_field_type_26_is_repeated,
  output [4:0]  io_out_bits_class_meta_field_type_26_field_type,
  output [15:0] io_out_bits_class_meta_field_type_26_sub_class_id,
  output        io_out_bits_class_meta_field_type_27_is_repeated,
  output [4:0]  io_out_bits_class_meta_field_type_27_field_type,
  output [15:0] io_out_bits_class_meta_field_type_27_sub_class_id,
  output        io_out_bits_class_meta_field_type_28_is_repeated,
  output [4:0]  io_out_bits_class_meta_field_type_28_field_type,
  output [15:0] io_out_bits_class_meta_field_type_28_sub_class_id,
  output        io_out_bits_class_meta_field_type_29_is_repeated,
  output [4:0]  io_out_bits_class_meta_field_type_29_field_type,
  output [15:0] io_out_bits_class_meta_field_type_29_sub_class_id,
  output        io_out_bits_class_meta_field_type_30_is_repeated,
  output [4:0]  io_out_bits_class_meta_field_type_30_field_type,
  output [15:0] io_out_bits_class_meta_field_type_30_sub_class_id,
  output        io_out_bits_class_meta_field_type_31_is_repeated,
  output [4:0]  io_out_bits_class_meta_field_type_31_field_type,
  output [15:0] io_out_bits_class_meta_field_type_31_sub_class_id,
  output        io_out_bits_class_meta_field_type_32_is_repeated,
  output [4:0]  io_out_bits_class_meta_field_type_32_field_type,
  output [15:0] io_out_bits_class_meta_field_type_32_sub_class_id
);
  wire  q_clock; // @[XQueue.scala 85:39]
  wire  q_reset; // @[XQueue.scala 85:39]
  wire  q_io_enq_ready; // @[XQueue.scala 85:39]
  wire  q_io_enq_valid; // @[XQueue.scala 85:39]
  wire [7:0] q_io_enq_bits_class_meta_max_field_num; // @[XQueue.scala 85:39]
  wire  q_io_enq_bits_class_meta_field_type_0_is_repeated; // @[XQueue.scala 85:39]
  wire [4:0] q_io_enq_bits_class_meta_field_type_0_field_type; // @[XQueue.scala 85:39]
  wire [15:0] q_io_enq_bits_class_meta_field_type_0_sub_class_id; // @[XQueue.scala 85:39]
  wire  q_io_enq_bits_class_meta_field_type_1_is_repeated; // @[XQueue.scala 85:39]
  wire [4:0] q_io_enq_bits_class_meta_field_type_1_field_type; // @[XQueue.scala 85:39]
  wire [15:0] q_io_enq_bits_class_meta_field_type_1_sub_class_id; // @[XQueue.scala 85:39]
  wire  q_io_enq_bits_class_meta_field_type_2_is_repeated; // @[XQueue.scala 85:39]
  wire [4:0] q_io_enq_bits_class_meta_field_type_2_field_type; // @[XQueue.scala 85:39]
  wire [15:0] q_io_enq_bits_class_meta_field_type_2_sub_class_id; // @[XQueue.scala 85:39]
  wire  q_io_enq_bits_class_meta_field_type_3_is_repeated; // @[XQueue.scala 85:39]
  wire [4:0] q_io_enq_bits_class_meta_field_type_3_field_type; // @[XQueue.scala 85:39]
  wire [15:0] q_io_enq_bits_class_meta_field_type_3_sub_class_id; // @[XQueue.scala 85:39]
  wire  q_io_enq_bits_class_meta_field_type_4_is_repeated; // @[XQueue.scala 85:39]
  wire [4:0] q_io_enq_bits_class_meta_field_type_4_field_type; // @[XQueue.scala 85:39]
  wire [15:0] q_io_enq_bits_class_meta_field_type_4_sub_class_id; // @[XQueue.scala 85:39]
  wire  q_io_enq_bits_class_meta_field_type_5_is_repeated; // @[XQueue.scala 85:39]
  wire [4:0] q_io_enq_bits_class_meta_field_type_5_field_type; // @[XQueue.scala 85:39]
  wire [15:0] q_io_enq_bits_class_meta_field_type_5_sub_class_id; // @[XQueue.scala 85:39]
  wire  q_io_enq_bits_class_meta_field_type_6_is_repeated; // @[XQueue.scala 85:39]
  wire [4:0] q_io_enq_bits_class_meta_field_type_6_field_type; // @[XQueue.scala 85:39]
  wire [15:0] q_io_enq_bits_class_meta_field_type_6_sub_class_id; // @[XQueue.scala 85:39]
  wire  q_io_enq_bits_class_meta_field_type_7_is_repeated; // @[XQueue.scala 85:39]
  wire [4:0] q_io_enq_bits_class_meta_field_type_7_field_type; // @[XQueue.scala 85:39]
  wire [15:0] q_io_enq_bits_class_meta_field_type_7_sub_class_id; // @[XQueue.scala 85:39]
  wire  q_io_enq_bits_class_meta_field_type_8_is_repeated; // @[XQueue.scala 85:39]
  wire [4:0] q_io_enq_bits_class_meta_field_type_8_field_type; // @[XQueue.scala 85:39]
  wire [15:0] q_io_enq_bits_class_meta_field_type_8_sub_class_id; // @[XQueue.scala 85:39]
  wire  q_io_enq_bits_class_meta_field_type_9_is_repeated; // @[XQueue.scala 85:39]
  wire [4:0] q_io_enq_bits_class_meta_field_type_9_field_type; // @[XQueue.scala 85:39]
  wire [15:0] q_io_enq_bits_class_meta_field_type_9_sub_class_id; // @[XQueue.scala 85:39]
  wire  q_io_enq_bits_class_meta_field_type_10_is_repeated; // @[XQueue.scala 85:39]
  wire [4:0] q_io_enq_bits_class_meta_field_type_10_field_type; // @[XQueue.scala 85:39]
  wire [15:0] q_io_enq_bits_class_meta_field_type_10_sub_class_id; // @[XQueue.scala 85:39]
  wire  q_io_enq_bits_class_meta_field_type_11_is_repeated; // @[XQueue.scala 85:39]
  wire [4:0] q_io_enq_bits_class_meta_field_type_11_field_type; // @[XQueue.scala 85:39]
  wire [15:0] q_io_enq_bits_class_meta_field_type_11_sub_class_id; // @[XQueue.scala 85:39]
  wire  q_io_enq_bits_class_meta_field_type_12_is_repeated; // @[XQueue.scala 85:39]
  wire [4:0] q_io_enq_bits_class_meta_field_type_12_field_type; // @[XQueue.scala 85:39]
  wire [15:0] q_io_enq_bits_class_meta_field_type_12_sub_class_id; // @[XQueue.scala 85:39]
  wire  q_io_enq_bits_class_meta_field_type_13_is_repeated; // @[XQueue.scala 85:39]
  wire [4:0] q_io_enq_bits_class_meta_field_type_13_field_type; // @[XQueue.scala 85:39]
  wire [15:0] q_io_enq_bits_class_meta_field_type_13_sub_class_id; // @[XQueue.scala 85:39]
  wire  q_io_enq_bits_class_meta_field_type_14_is_repeated; // @[XQueue.scala 85:39]
  wire [4:0] q_io_enq_bits_class_meta_field_type_14_field_type; // @[XQueue.scala 85:39]
  wire [15:0] q_io_enq_bits_class_meta_field_type_14_sub_class_id; // @[XQueue.scala 85:39]
  wire  q_io_enq_bits_class_meta_field_type_15_is_repeated; // @[XQueue.scala 85:39]
  wire [4:0] q_io_enq_bits_class_meta_field_type_15_field_type; // @[XQueue.scala 85:39]
  wire [15:0] q_io_enq_bits_class_meta_field_type_15_sub_class_id; // @[XQueue.scala 85:39]
  wire  q_io_enq_bits_class_meta_field_type_16_is_repeated; // @[XQueue.scala 85:39]
  wire [4:0] q_io_enq_bits_class_meta_field_type_16_field_type; // @[XQueue.scala 85:39]
  wire [15:0] q_io_enq_bits_class_meta_field_type_16_sub_class_id; // @[XQueue.scala 85:39]
  wire  q_io_enq_bits_class_meta_field_type_17_is_repeated; // @[XQueue.scala 85:39]
  wire [4:0] q_io_enq_bits_class_meta_field_type_17_field_type; // @[XQueue.scala 85:39]
  wire [15:0] q_io_enq_bits_class_meta_field_type_17_sub_class_id; // @[XQueue.scala 85:39]
  wire  q_io_enq_bits_class_meta_field_type_18_is_repeated; // @[XQueue.scala 85:39]
  wire [4:0] q_io_enq_bits_class_meta_field_type_18_field_type; // @[XQueue.scala 85:39]
  wire [15:0] q_io_enq_bits_class_meta_field_type_18_sub_class_id; // @[XQueue.scala 85:39]
  wire  q_io_enq_bits_class_meta_field_type_19_is_repeated; // @[XQueue.scala 85:39]
  wire [4:0] q_io_enq_bits_class_meta_field_type_19_field_type; // @[XQueue.scala 85:39]
  wire [15:0] q_io_enq_bits_class_meta_field_type_19_sub_class_id; // @[XQueue.scala 85:39]
  wire  q_io_enq_bits_class_meta_field_type_20_is_repeated; // @[XQueue.scala 85:39]
  wire [4:0] q_io_enq_bits_class_meta_field_type_20_field_type; // @[XQueue.scala 85:39]
  wire [15:0] q_io_enq_bits_class_meta_field_type_20_sub_class_id; // @[XQueue.scala 85:39]
  wire  q_io_enq_bits_class_meta_field_type_21_is_repeated; // @[XQueue.scala 85:39]
  wire [4:0] q_io_enq_bits_class_meta_field_type_21_field_type; // @[XQueue.scala 85:39]
  wire [15:0] q_io_enq_bits_class_meta_field_type_21_sub_class_id; // @[XQueue.scala 85:39]
  wire  q_io_enq_bits_class_meta_field_type_22_is_repeated; // @[XQueue.scala 85:39]
  wire [4:0] q_io_enq_bits_class_meta_field_type_22_field_type; // @[XQueue.scala 85:39]
  wire [15:0] q_io_enq_bits_class_meta_field_type_22_sub_class_id; // @[XQueue.scala 85:39]
  wire  q_io_enq_bits_class_meta_field_type_23_is_repeated; // @[XQueue.scala 85:39]
  wire [4:0] q_io_enq_bits_class_meta_field_type_23_field_type; // @[XQueue.scala 85:39]
  wire [15:0] q_io_enq_bits_class_meta_field_type_23_sub_class_id; // @[XQueue.scala 85:39]
  wire  q_io_enq_bits_class_meta_field_type_24_is_repeated; // @[XQueue.scala 85:39]
  wire [4:0] q_io_enq_bits_class_meta_field_type_24_field_type; // @[XQueue.scala 85:39]
  wire [15:0] q_io_enq_bits_class_meta_field_type_24_sub_class_id; // @[XQueue.scala 85:39]
  wire  q_io_enq_bits_class_meta_field_type_25_is_repeated; // @[XQueue.scala 85:39]
  wire [4:0] q_io_enq_bits_class_meta_field_type_25_field_type; // @[XQueue.scala 85:39]
  wire [15:0] q_io_enq_bits_class_meta_field_type_25_sub_class_id; // @[XQueue.scala 85:39]
  wire  q_io_enq_bits_class_meta_field_type_26_is_repeated; // @[XQueue.scala 85:39]
  wire [4:0] q_io_enq_bits_class_meta_field_type_26_field_type; // @[XQueue.scala 85:39]
  wire [15:0] q_io_enq_bits_class_meta_field_type_26_sub_class_id; // @[XQueue.scala 85:39]
  wire  q_io_enq_bits_class_meta_field_type_27_is_repeated; // @[XQueue.scala 85:39]
  wire [4:0] q_io_enq_bits_class_meta_field_type_27_field_type; // @[XQueue.scala 85:39]
  wire [15:0] q_io_enq_bits_class_meta_field_type_27_sub_class_id; // @[XQueue.scala 85:39]
  wire  q_io_enq_bits_class_meta_field_type_28_is_repeated; // @[XQueue.scala 85:39]
  wire [4:0] q_io_enq_bits_class_meta_field_type_28_field_type; // @[XQueue.scala 85:39]
  wire [15:0] q_io_enq_bits_class_meta_field_type_28_sub_class_id; // @[XQueue.scala 85:39]
  wire  q_io_enq_bits_class_meta_field_type_29_is_repeated; // @[XQueue.scala 85:39]
  wire [4:0] q_io_enq_bits_class_meta_field_type_29_field_type; // @[XQueue.scala 85:39]
  wire [15:0] q_io_enq_bits_class_meta_field_type_29_sub_class_id; // @[XQueue.scala 85:39]
  wire  q_io_enq_bits_class_meta_field_type_30_is_repeated; // @[XQueue.scala 85:39]
  wire [4:0] q_io_enq_bits_class_meta_field_type_30_field_type; // @[XQueue.scala 85:39]
  wire [15:0] q_io_enq_bits_class_meta_field_type_30_sub_class_id; // @[XQueue.scala 85:39]
  wire  q_io_enq_bits_class_meta_field_type_31_is_repeated; // @[XQueue.scala 85:39]
  wire [4:0] q_io_enq_bits_class_meta_field_type_31_field_type; // @[XQueue.scala 85:39]
  wire [15:0] q_io_enq_bits_class_meta_field_type_31_sub_class_id; // @[XQueue.scala 85:39]
  wire  q_io_enq_bits_class_meta_field_type_32_is_repeated; // @[XQueue.scala 85:39]
  wire [4:0] q_io_enq_bits_class_meta_field_type_32_field_type; // @[XQueue.scala 85:39]
  wire [15:0] q_io_enq_bits_class_meta_field_type_32_sub_class_id; // @[XQueue.scala 85:39]
  wire  q_io_deq_ready; // @[XQueue.scala 85:39]
  wire  q_io_deq_valid; // @[XQueue.scala 85:39]
  wire [7:0] q_io_deq_bits_class_meta_max_field_num; // @[XQueue.scala 85:39]
  wire  q_io_deq_bits_class_meta_field_type_0_is_repeated; // @[XQueue.scala 85:39]
  wire [4:0] q_io_deq_bits_class_meta_field_type_0_field_type; // @[XQueue.scala 85:39]
  wire [15:0] q_io_deq_bits_class_meta_field_type_0_sub_class_id; // @[XQueue.scala 85:39]
  wire  q_io_deq_bits_class_meta_field_type_1_is_repeated; // @[XQueue.scala 85:39]
  wire [4:0] q_io_deq_bits_class_meta_field_type_1_field_type; // @[XQueue.scala 85:39]
  wire [15:0] q_io_deq_bits_class_meta_field_type_1_sub_class_id; // @[XQueue.scala 85:39]
  wire  q_io_deq_bits_class_meta_field_type_2_is_repeated; // @[XQueue.scala 85:39]
  wire [4:0] q_io_deq_bits_class_meta_field_type_2_field_type; // @[XQueue.scala 85:39]
  wire [15:0] q_io_deq_bits_class_meta_field_type_2_sub_class_id; // @[XQueue.scala 85:39]
  wire  q_io_deq_bits_class_meta_field_type_3_is_repeated; // @[XQueue.scala 85:39]
  wire [4:0] q_io_deq_bits_class_meta_field_type_3_field_type; // @[XQueue.scala 85:39]
  wire [15:0] q_io_deq_bits_class_meta_field_type_3_sub_class_id; // @[XQueue.scala 85:39]
  wire  q_io_deq_bits_class_meta_field_type_4_is_repeated; // @[XQueue.scala 85:39]
  wire [4:0] q_io_deq_bits_class_meta_field_type_4_field_type; // @[XQueue.scala 85:39]
  wire [15:0] q_io_deq_bits_class_meta_field_type_4_sub_class_id; // @[XQueue.scala 85:39]
  wire  q_io_deq_bits_class_meta_field_type_5_is_repeated; // @[XQueue.scala 85:39]
  wire [4:0] q_io_deq_bits_class_meta_field_type_5_field_type; // @[XQueue.scala 85:39]
  wire [15:0] q_io_deq_bits_class_meta_field_type_5_sub_class_id; // @[XQueue.scala 85:39]
  wire  q_io_deq_bits_class_meta_field_type_6_is_repeated; // @[XQueue.scala 85:39]
  wire [4:0] q_io_deq_bits_class_meta_field_type_6_field_type; // @[XQueue.scala 85:39]
  wire [15:0] q_io_deq_bits_class_meta_field_type_6_sub_class_id; // @[XQueue.scala 85:39]
  wire  q_io_deq_bits_class_meta_field_type_7_is_repeated; // @[XQueue.scala 85:39]
  wire [4:0] q_io_deq_bits_class_meta_field_type_7_field_type; // @[XQueue.scala 85:39]
  wire [15:0] q_io_deq_bits_class_meta_field_type_7_sub_class_id; // @[XQueue.scala 85:39]
  wire  q_io_deq_bits_class_meta_field_type_8_is_repeated; // @[XQueue.scala 85:39]
  wire [4:0] q_io_deq_bits_class_meta_field_type_8_field_type; // @[XQueue.scala 85:39]
  wire [15:0] q_io_deq_bits_class_meta_field_type_8_sub_class_id; // @[XQueue.scala 85:39]
  wire  q_io_deq_bits_class_meta_field_type_9_is_repeated; // @[XQueue.scala 85:39]
  wire [4:0] q_io_deq_bits_class_meta_field_type_9_field_type; // @[XQueue.scala 85:39]
  wire [15:0] q_io_deq_bits_class_meta_field_type_9_sub_class_id; // @[XQueue.scala 85:39]
  wire  q_io_deq_bits_class_meta_field_type_10_is_repeated; // @[XQueue.scala 85:39]
  wire [4:0] q_io_deq_bits_class_meta_field_type_10_field_type; // @[XQueue.scala 85:39]
  wire [15:0] q_io_deq_bits_class_meta_field_type_10_sub_class_id; // @[XQueue.scala 85:39]
  wire  q_io_deq_bits_class_meta_field_type_11_is_repeated; // @[XQueue.scala 85:39]
  wire [4:0] q_io_deq_bits_class_meta_field_type_11_field_type; // @[XQueue.scala 85:39]
  wire [15:0] q_io_deq_bits_class_meta_field_type_11_sub_class_id; // @[XQueue.scala 85:39]
  wire  q_io_deq_bits_class_meta_field_type_12_is_repeated; // @[XQueue.scala 85:39]
  wire [4:0] q_io_deq_bits_class_meta_field_type_12_field_type; // @[XQueue.scala 85:39]
  wire [15:0] q_io_deq_bits_class_meta_field_type_12_sub_class_id; // @[XQueue.scala 85:39]
  wire  q_io_deq_bits_class_meta_field_type_13_is_repeated; // @[XQueue.scala 85:39]
  wire [4:0] q_io_deq_bits_class_meta_field_type_13_field_type; // @[XQueue.scala 85:39]
  wire [15:0] q_io_deq_bits_class_meta_field_type_13_sub_class_id; // @[XQueue.scala 85:39]
  wire  q_io_deq_bits_class_meta_field_type_14_is_repeated; // @[XQueue.scala 85:39]
  wire [4:0] q_io_deq_bits_class_meta_field_type_14_field_type; // @[XQueue.scala 85:39]
  wire [15:0] q_io_deq_bits_class_meta_field_type_14_sub_class_id; // @[XQueue.scala 85:39]
  wire  q_io_deq_bits_class_meta_field_type_15_is_repeated; // @[XQueue.scala 85:39]
  wire [4:0] q_io_deq_bits_class_meta_field_type_15_field_type; // @[XQueue.scala 85:39]
  wire [15:0] q_io_deq_bits_class_meta_field_type_15_sub_class_id; // @[XQueue.scala 85:39]
  wire  q_io_deq_bits_class_meta_field_type_16_is_repeated; // @[XQueue.scala 85:39]
  wire [4:0] q_io_deq_bits_class_meta_field_type_16_field_type; // @[XQueue.scala 85:39]
  wire [15:0] q_io_deq_bits_class_meta_field_type_16_sub_class_id; // @[XQueue.scala 85:39]
  wire  q_io_deq_bits_class_meta_field_type_17_is_repeated; // @[XQueue.scala 85:39]
  wire [4:0] q_io_deq_bits_class_meta_field_type_17_field_type; // @[XQueue.scala 85:39]
  wire [15:0] q_io_deq_bits_class_meta_field_type_17_sub_class_id; // @[XQueue.scala 85:39]
  wire  q_io_deq_bits_class_meta_field_type_18_is_repeated; // @[XQueue.scala 85:39]
  wire [4:0] q_io_deq_bits_class_meta_field_type_18_field_type; // @[XQueue.scala 85:39]
  wire [15:0] q_io_deq_bits_class_meta_field_type_18_sub_class_id; // @[XQueue.scala 85:39]
  wire  q_io_deq_bits_class_meta_field_type_19_is_repeated; // @[XQueue.scala 85:39]
  wire [4:0] q_io_deq_bits_class_meta_field_type_19_field_type; // @[XQueue.scala 85:39]
  wire [15:0] q_io_deq_bits_class_meta_field_type_19_sub_class_id; // @[XQueue.scala 85:39]
  wire  q_io_deq_bits_class_meta_field_type_20_is_repeated; // @[XQueue.scala 85:39]
  wire [4:0] q_io_deq_bits_class_meta_field_type_20_field_type; // @[XQueue.scala 85:39]
  wire [15:0] q_io_deq_bits_class_meta_field_type_20_sub_class_id; // @[XQueue.scala 85:39]
  wire  q_io_deq_bits_class_meta_field_type_21_is_repeated; // @[XQueue.scala 85:39]
  wire [4:0] q_io_deq_bits_class_meta_field_type_21_field_type; // @[XQueue.scala 85:39]
  wire [15:0] q_io_deq_bits_class_meta_field_type_21_sub_class_id; // @[XQueue.scala 85:39]
  wire  q_io_deq_bits_class_meta_field_type_22_is_repeated; // @[XQueue.scala 85:39]
  wire [4:0] q_io_deq_bits_class_meta_field_type_22_field_type; // @[XQueue.scala 85:39]
  wire [15:0] q_io_deq_bits_class_meta_field_type_22_sub_class_id; // @[XQueue.scala 85:39]
  wire  q_io_deq_bits_class_meta_field_type_23_is_repeated; // @[XQueue.scala 85:39]
  wire [4:0] q_io_deq_bits_class_meta_field_type_23_field_type; // @[XQueue.scala 85:39]
  wire [15:0] q_io_deq_bits_class_meta_field_type_23_sub_class_id; // @[XQueue.scala 85:39]
  wire  q_io_deq_bits_class_meta_field_type_24_is_repeated; // @[XQueue.scala 85:39]
  wire [4:0] q_io_deq_bits_class_meta_field_type_24_field_type; // @[XQueue.scala 85:39]
  wire [15:0] q_io_deq_bits_class_meta_field_type_24_sub_class_id; // @[XQueue.scala 85:39]
  wire  q_io_deq_bits_class_meta_field_type_25_is_repeated; // @[XQueue.scala 85:39]
  wire [4:0] q_io_deq_bits_class_meta_field_type_25_field_type; // @[XQueue.scala 85:39]
  wire [15:0] q_io_deq_bits_class_meta_field_type_25_sub_class_id; // @[XQueue.scala 85:39]
  wire  q_io_deq_bits_class_meta_field_type_26_is_repeated; // @[XQueue.scala 85:39]
  wire [4:0] q_io_deq_bits_class_meta_field_type_26_field_type; // @[XQueue.scala 85:39]
  wire [15:0] q_io_deq_bits_class_meta_field_type_26_sub_class_id; // @[XQueue.scala 85:39]
  wire  q_io_deq_bits_class_meta_field_type_27_is_repeated; // @[XQueue.scala 85:39]
  wire [4:0] q_io_deq_bits_class_meta_field_type_27_field_type; // @[XQueue.scala 85:39]
  wire [15:0] q_io_deq_bits_class_meta_field_type_27_sub_class_id; // @[XQueue.scala 85:39]
  wire  q_io_deq_bits_class_meta_field_type_28_is_repeated; // @[XQueue.scala 85:39]
  wire [4:0] q_io_deq_bits_class_meta_field_type_28_field_type; // @[XQueue.scala 85:39]
  wire [15:0] q_io_deq_bits_class_meta_field_type_28_sub_class_id; // @[XQueue.scala 85:39]
  wire  q_io_deq_bits_class_meta_field_type_29_is_repeated; // @[XQueue.scala 85:39]
  wire [4:0] q_io_deq_bits_class_meta_field_type_29_field_type; // @[XQueue.scala 85:39]
  wire [15:0] q_io_deq_bits_class_meta_field_type_29_sub_class_id; // @[XQueue.scala 85:39]
  wire  q_io_deq_bits_class_meta_field_type_30_is_repeated; // @[XQueue.scala 85:39]
  wire [4:0] q_io_deq_bits_class_meta_field_type_30_field_type; // @[XQueue.scala 85:39]
  wire [15:0] q_io_deq_bits_class_meta_field_type_30_sub_class_id; // @[XQueue.scala 85:39]
  wire  q_io_deq_bits_class_meta_field_type_31_is_repeated; // @[XQueue.scala 85:39]
  wire [4:0] q_io_deq_bits_class_meta_field_type_31_field_type; // @[XQueue.scala 85:39]
  wire [15:0] q_io_deq_bits_class_meta_field_type_31_sub_class_id; // @[XQueue.scala 85:39]
  wire  q_io_deq_bits_class_meta_field_type_32_is_repeated; // @[XQueue.scala 85:39]
  wire [4:0] q_io_deq_bits_class_meta_field_type_32_field_type; // @[XQueue.scala 85:39]
  wire [15:0] q_io_deq_bits_class_meta_field_type_32_sub_class_id; // @[XQueue.scala 85:39]
  Queue_5 q ( // @[XQueue.scala 85:39]
    .clock(q_clock),
    .reset(q_reset),
    .io_enq_ready(q_io_enq_ready),
    .io_enq_valid(q_io_enq_valid),
    .io_enq_bits_class_meta_max_field_num(q_io_enq_bits_class_meta_max_field_num),
    .io_enq_bits_class_meta_field_type_0_is_repeated(q_io_enq_bits_class_meta_field_type_0_is_repeated),
    .io_enq_bits_class_meta_field_type_0_field_type(q_io_enq_bits_class_meta_field_type_0_field_type),
    .io_enq_bits_class_meta_field_type_0_sub_class_id(q_io_enq_bits_class_meta_field_type_0_sub_class_id),
    .io_enq_bits_class_meta_field_type_1_is_repeated(q_io_enq_bits_class_meta_field_type_1_is_repeated),
    .io_enq_bits_class_meta_field_type_1_field_type(q_io_enq_bits_class_meta_field_type_1_field_type),
    .io_enq_bits_class_meta_field_type_1_sub_class_id(q_io_enq_bits_class_meta_field_type_1_sub_class_id),
    .io_enq_bits_class_meta_field_type_2_is_repeated(q_io_enq_bits_class_meta_field_type_2_is_repeated),
    .io_enq_bits_class_meta_field_type_2_field_type(q_io_enq_bits_class_meta_field_type_2_field_type),
    .io_enq_bits_class_meta_field_type_2_sub_class_id(q_io_enq_bits_class_meta_field_type_2_sub_class_id),
    .io_enq_bits_class_meta_field_type_3_is_repeated(q_io_enq_bits_class_meta_field_type_3_is_repeated),
    .io_enq_bits_class_meta_field_type_3_field_type(q_io_enq_bits_class_meta_field_type_3_field_type),
    .io_enq_bits_class_meta_field_type_3_sub_class_id(q_io_enq_bits_class_meta_field_type_3_sub_class_id),
    .io_enq_bits_class_meta_field_type_4_is_repeated(q_io_enq_bits_class_meta_field_type_4_is_repeated),
    .io_enq_bits_class_meta_field_type_4_field_type(q_io_enq_bits_class_meta_field_type_4_field_type),
    .io_enq_bits_class_meta_field_type_4_sub_class_id(q_io_enq_bits_class_meta_field_type_4_sub_class_id),
    .io_enq_bits_class_meta_field_type_5_is_repeated(q_io_enq_bits_class_meta_field_type_5_is_repeated),
    .io_enq_bits_class_meta_field_type_5_field_type(q_io_enq_bits_class_meta_field_type_5_field_type),
    .io_enq_bits_class_meta_field_type_5_sub_class_id(q_io_enq_bits_class_meta_field_type_5_sub_class_id),
    .io_enq_bits_class_meta_field_type_6_is_repeated(q_io_enq_bits_class_meta_field_type_6_is_repeated),
    .io_enq_bits_class_meta_field_type_6_field_type(q_io_enq_bits_class_meta_field_type_6_field_type),
    .io_enq_bits_class_meta_field_type_6_sub_class_id(q_io_enq_bits_class_meta_field_type_6_sub_class_id),
    .io_enq_bits_class_meta_field_type_7_is_repeated(q_io_enq_bits_class_meta_field_type_7_is_repeated),
    .io_enq_bits_class_meta_field_type_7_field_type(q_io_enq_bits_class_meta_field_type_7_field_type),
    .io_enq_bits_class_meta_field_type_7_sub_class_id(q_io_enq_bits_class_meta_field_type_7_sub_class_id),
    .io_enq_bits_class_meta_field_type_8_is_repeated(q_io_enq_bits_class_meta_field_type_8_is_repeated),
    .io_enq_bits_class_meta_field_type_8_field_type(q_io_enq_bits_class_meta_field_type_8_field_type),
    .io_enq_bits_class_meta_field_type_8_sub_class_id(q_io_enq_bits_class_meta_field_type_8_sub_class_id),
    .io_enq_bits_class_meta_field_type_9_is_repeated(q_io_enq_bits_class_meta_field_type_9_is_repeated),
    .io_enq_bits_class_meta_field_type_9_field_type(q_io_enq_bits_class_meta_field_type_9_field_type),
    .io_enq_bits_class_meta_field_type_9_sub_class_id(q_io_enq_bits_class_meta_field_type_9_sub_class_id),
    .io_enq_bits_class_meta_field_type_10_is_repeated(q_io_enq_bits_class_meta_field_type_10_is_repeated),
    .io_enq_bits_class_meta_field_type_10_field_type(q_io_enq_bits_class_meta_field_type_10_field_type),
    .io_enq_bits_class_meta_field_type_10_sub_class_id(q_io_enq_bits_class_meta_field_type_10_sub_class_id),
    .io_enq_bits_class_meta_field_type_11_is_repeated(q_io_enq_bits_class_meta_field_type_11_is_repeated),
    .io_enq_bits_class_meta_field_type_11_field_type(q_io_enq_bits_class_meta_field_type_11_field_type),
    .io_enq_bits_class_meta_field_type_11_sub_class_id(q_io_enq_bits_class_meta_field_type_11_sub_class_id),
    .io_enq_bits_class_meta_field_type_12_is_repeated(q_io_enq_bits_class_meta_field_type_12_is_repeated),
    .io_enq_bits_class_meta_field_type_12_field_type(q_io_enq_bits_class_meta_field_type_12_field_type),
    .io_enq_bits_class_meta_field_type_12_sub_class_id(q_io_enq_bits_class_meta_field_type_12_sub_class_id),
    .io_enq_bits_class_meta_field_type_13_is_repeated(q_io_enq_bits_class_meta_field_type_13_is_repeated),
    .io_enq_bits_class_meta_field_type_13_field_type(q_io_enq_bits_class_meta_field_type_13_field_type),
    .io_enq_bits_class_meta_field_type_13_sub_class_id(q_io_enq_bits_class_meta_field_type_13_sub_class_id),
    .io_enq_bits_class_meta_field_type_14_is_repeated(q_io_enq_bits_class_meta_field_type_14_is_repeated),
    .io_enq_bits_class_meta_field_type_14_field_type(q_io_enq_bits_class_meta_field_type_14_field_type),
    .io_enq_bits_class_meta_field_type_14_sub_class_id(q_io_enq_bits_class_meta_field_type_14_sub_class_id),
    .io_enq_bits_class_meta_field_type_15_is_repeated(q_io_enq_bits_class_meta_field_type_15_is_repeated),
    .io_enq_bits_class_meta_field_type_15_field_type(q_io_enq_bits_class_meta_field_type_15_field_type),
    .io_enq_bits_class_meta_field_type_15_sub_class_id(q_io_enq_bits_class_meta_field_type_15_sub_class_id),
    .io_enq_bits_class_meta_field_type_16_is_repeated(q_io_enq_bits_class_meta_field_type_16_is_repeated),
    .io_enq_bits_class_meta_field_type_16_field_type(q_io_enq_bits_class_meta_field_type_16_field_type),
    .io_enq_bits_class_meta_field_type_16_sub_class_id(q_io_enq_bits_class_meta_field_type_16_sub_class_id),
    .io_enq_bits_class_meta_field_type_17_is_repeated(q_io_enq_bits_class_meta_field_type_17_is_repeated),
    .io_enq_bits_class_meta_field_type_17_field_type(q_io_enq_bits_class_meta_field_type_17_field_type),
    .io_enq_bits_class_meta_field_type_17_sub_class_id(q_io_enq_bits_class_meta_field_type_17_sub_class_id),
    .io_enq_bits_class_meta_field_type_18_is_repeated(q_io_enq_bits_class_meta_field_type_18_is_repeated),
    .io_enq_bits_class_meta_field_type_18_field_type(q_io_enq_bits_class_meta_field_type_18_field_type),
    .io_enq_bits_class_meta_field_type_18_sub_class_id(q_io_enq_bits_class_meta_field_type_18_sub_class_id),
    .io_enq_bits_class_meta_field_type_19_is_repeated(q_io_enq_bits_class_meta_field_type_19_is_repeated),
    .io_enq_bits_class_meta_field_type_19_field_type(q_io_enq_bits_class_meta_field_type_19_field_type),
    .io_enq_bits_class_meta_field_type_19_sub_class_id(q_io_enq_bits_class_meta_field_type_19_sub_class_id),
    .io_enq_bits_class_meta_field_type_20_is_repeated(q_io_enq_bits_class_meta_field_type_20_is_repeated),
    .io_enq_bits_class_meta_field_type_20_field_type(q_io_enq_bits_class_meta_field_type_20_field_type),
    .io_enq_bits_class_meta_field_type_20_sub_class_id(q_io_enq_bits_class_meta_field_type_20_sub_class_id),
    .io_enq_bits_class_meta_field_type_21_is_repeated(q_io_enq_bits_class_meta_field_type_21_is_repeated),
    .io_enq_bits_class_meta_field_type_21_field_type(q_io_enq_bits_class_meta_field_type_21_field_type),
    .io_enq_bits_class_meta_field_type_21_sub_class_id(q_io_enq_bits_class_meta_field_type_21_sub_class_id),
    .io_enq_bits_class_meta_field_type_22_is_repeated(q_io_enq_bits_class_meta_field_type_22_is_repeated),
    .io_enq_bits_class_meta_field_type_22_field_type(q_io_enq_bits_class_meta_field_type_22_field_type),
    .io_enq_bits_class_meta_field_type_22_sub_class_id(q_io_enq_bits_class_meta_field_type_22_sub_class_id),
    .io_enq_bits_class_meta_field_type_23_is_repeated(q_io_enq_bits_class_meta_field_type_23_is_repeated),
    .io_enq_bits_class_meta_field_type_23_field_type(q_io_enq_bits_class_meta_field_type_23_field_type),
    .io_enq_bits_class_meta_field_type_23_sub_class_id(q_io_enq_bits_class_meta_field_type_23_sub_class_id),
    .io_enq_bits_class_meta_field_type_24_is_repeated(q_io_enq_bits_class_meta_field_type_24_is_repeated),
    .io_enq_bits_class_meta_field_type_24_field_type(q_io_enq_bits_class_meta_field_type_24_field_type),
    .io_enq_bits_class_meta_field_type_24_sub_class_id(q_io_enq_bits_class_meta_field_type_24_sub_class_id),
    .io_enq_bits_class_meta_field_type_25_is_repeated(q_io_enq_bits_class_meta_field_type_25_is_repeated),
    .io_enq_bits_class_meta_field_type_25_field_type(q_io_enq_bits_class_meta_field_type_25_field_type),
    .io_enq_bits_class_meta_field_type_25_sub_class_id(q_io_enq_bits_class_meta_field_type_25_sub_class_id),
    .io_enq_bits_class_meta_field_type_26_is_repeated(q_io_enq_bits_class_meta_field_type_26_is_repeated),
    .io_enq_bits_class_meta_field_type_26_field_type(q_io_enq_bits_class_meta_field_type_26_field_type),
    .io_enq_bits_class_meta_field_type_26_sub_class_id(q_io_enq_bits_class_meta_field_type_26_sub_class_id),
    .io_enq_bits_class_meta_field_type_27_is_repeated(q_io_enq_bits_class_meta_field_type_27_is_repeated),
    .io_enq_bits_class_meta_field_type_27_field_type(q_io_enq_bits_class_meta_field_type_27_field_type),
    .io_enq_bits_class_meta_field_type_27_sub_class_id(q_io_enq_bits_class_meta_field_type_27_sub_class_id),
    .io_enq_bits_class_meta_field_type_28_is_repeated(q_io_enq_bits_class_meta_field_type_28_is_repeated),
    .io_enq_bits_class_meta_field_type_28_field_type(q_io_enq_bits_class_meta_field_type_28_field_type),
    .io_enq_bits_class_meta_field_type_28_sub_class_id(q_io_enq_bits_class_meta_field_type_28_sub_class_id),
    .io_enq_bits_class_meta_field_type_29_is_repeated(q_io_enq_bits_class_meta_field_type_29_is_repeated),
    .io_enq_bits_class_meta_field_type_29_field_type(q_io_enq_bits_class_meta_field_type_29_field_type),
    .io_enq_bits_class_meta_field_type_29_sub_class_id(q_io_enq_bits_class_meta_field_type_29_sub_class_id),
    .io_enq_bits_class_meta_field_type_30_is_repeated(q_io_enq_bits_class_meta_field_type_30_is_repeated),
    .io_enq_bits_class_meta_field_type_30_field_type(q_io_enq_bits_class_meta_field_type_30_field_type),
    .io_enq_bits_class_meta_field_type_30_sub_class_id(q_io_enq_bits_class_meta_field_type_30_sub_class_id),
    .io_enq_bits_class_meta_field_type_31_is_repeated(q_io_enq_bits_class_meta_field_type_31_is_repeated),
    .io_enq_bits_class_meta_field_type_31_field_type(q_io_enq_bits_class_meta_field_type_31_field_type),
    .io_enq_bits_class_meta_field_type_31_sub_class_id(q_io_enq_bits_class_meta_field_type_31_sub_class_id),
    .io_enq_bits_class_meta_field_type_32_is_repeated(q_io_enq_bits_class_meta_field_type_32_is_repeated),
    .io_enq_bits_class_meta_field_type_32_field_type(q_io_enq_bits_class_meta_field_type_32_field_type),
    .io_enq_bits_class_meta_field_type_32_sub_class_id(q_io_enq_bits_class_meta_field_type_32_sub_class_id),
    .io_deq_ready(q_io_deq_ready),
    .io_deq_valid(q_io_deq_valid),
    .io_deq_bits_class_meta_max_field_num(q_io_deq_bits_class_meta_max_field_num),
    .io_deq_bits_class_meta_field_type_0_is_repeated(q_io_deq_bits_class_meta_field_type_0_is_repeated),
    .io_deq_bits_class_meta_field_type_0_field_type(q_io_deq_bits_class_meta_field_type_0_field_type),
    .io_deq_bits_class_meta_field_type_0_sub_class_id(q_io_deq_bits_class_meta_field_type_0_sub_class_id),
    .io_deq_bits_class_meta_field_type_1_is_repeated(q_io_deq_bits_class_meta_field_type_1_is_repeated),
    .io_deq_bits_class_meta_field_type_1_field_type(q_io_deq_bits_class_meta_field_type_1_field_type),
    .io_deq_bits_class_meta_field_type_1_sub_class_id(q_io_deq_bits_class_meta_field_type_1_sub_class_id),
    .io_deq_bits_class_meta_field_type_2_is_repeated(q_io_deq_bits_class_meta_field_type_2_is_repeated),
    .io_deq_bits_class_meta_field_type_2_field_type(q_io_deq_bits_class_meta_field_type_2_field_type),
    .io_deq_bits_class_meta_field_type_2_sub_class_id(q_io_deq_bits_class_meta_field_type_2_sub_class_id),
    .io_deq_bits_class_meta_field_type_3_is_repeated(q_io_deq_bits_class_meta_field_type_3_is_repeated),
    .io_deq_bits_class_meta_field_type_3_field_type(q_io_deq_bits_class_meta_field_type_3_field_type),
    .io_deq_bits_class_meta_field_type_3_sub_class_id(q_io_deq_bits_class_meta_field_type_3_sub_class_id),
    .io_deq_bits_class_meta_field_type_4_is_repeated(q_io_deq_bits_class_meta_field_type_4_is_repeated),
    .io_deq_bits_class_meta_field_type_4_field_type(q_io_deq_bits_class_meta_field_type_4_field_type),
    .io_deq_bits_class_meta_field_type_4_sub_class_id(q_io_deq_bits_class_meta_field_type_4_sub_class_id),
    .io_deq_bits_class_meta_field_type_5_is_repeated(q_io_deq_bits_class_meta_field_type_5_is_repeated),
    .io_deq_bits_class_meta_field_type_5_field_type(q_io_deq_bits_class_meta_field_type_5_field_type),
    .io_deq_bits_class_meta_field_type_5_sub_class_id(q_io_deq_bits_class_meta_field_type_5_sub_class_id),
    .io_deq_bits_class_meta_field_type_6_is_repeated(q_io_deq_bits_class_meta_field_type_6_is_repeated),
    .io_deq_bits_class_meta_field_type_6_field_type(q_io_deq_bits_class_meta_field_type_6_field_type),
    .io_deq_bits_class_meta_field_type_6_sub_class_id(q_io_deq_bits_class_meta_field_type_6_sub_class_id),
    .io_deq_bits_class_meta_field_type_7_is_repeated(q_io_deq_bits_class_meta_field_type_7_is_repeated),
    .io_deq_bits_class_meta_field_type_7_field_type(q_io_deq_bits_class_meta_field_type_7_field_type),
    .io_deq_bits_class_meta_field_type_7_sub_class_id(q_io_deq_bits_class_meta_field_type_7_sub_class_id),
    .io_deq_bits_class_meta_field_type_8_is_repeated(q_io_deq_bits_class_meta_field_type_8_is_repeated),
    .io_deq_bits_class_meta_field_type_8_field_type(q_io_deq_bits_class_meta_field_type_8_field_type),
    .io_deq_bits_class_meta_field_type_8_sub_class_id(q_io_deq_bits_class_meta_field_type_8_sub_class_id),
    .io_deq_bits_class_meta_field_type_9_is_repeated(q_io_deq_bits_class_meta_field_type_9_is_repeated),
    .io_deq_bits_class_meta_field_type_9_field_type(q_io_deq_bits_class_meta_field_type_9_field_type),
    .io_deq_bits_class_meta_field_type_9_sub_class_id(q_io_deq_bits_class_meta_field_type_9_sub_class_id),
    .io_deq_bits_class_meta_field_type_10_is_repeated(q_io_deq_bits_class_meta_field_type_10_is_repeated),
    .io_deq_bits_class_meta_field_type_10_field_type(q_io_deq_bits_class_meta_field_type_10_field_type),
    .io_deq_bits_class_meta_field_type_10_sub_class_id(q_io_deq_bits_class_meta_field_type_10_sub_class_id),
    .io_deq_bits_class_meta_field_type_11_is_repeated(q_io_deq_bits_class_meta_field_type_11_is_repeated),
    .io_deq_bits_class_meta_field_type_11_field_type(q_io_deq_bits_class_meta_field_type_11_field_type),
    .io_deq_bits_class_meta_field_type_11_sub_class_id(q_io_deq_bits_class_meta_field_type_11_sub_class_id),
    .io_deq_bits_class_meta_field_type_12_is_repeated(q_io_deq_bits_class_meta_field_type_12_is_repeated),
    .io_deq_bits_class_meta_field_type_12_field_type(q_io_deq_bits_class_meta_field_type_12_field_type),
    .io_deq_bits_class_meta_field_type_12_sub_class_id(q_io_deq_bits_class_meta_field_type_12_sub_class_id),
    .io_deq_bits_class_meta_field_type_13_is_repeated(q_io_deq_bits_class_meta_field_type_13_is_repeated),
    .io_deq_bits_class_meta_field_type_13_field_type(q_io_deq_bits_class_meta_field_type_13_field_type),
    .io_deq_bits_class_meta_field_type_13_sub_class_id(q_io_deq_bits_class_meta_field_type_13_sub_class_id),
    .io_deq_bits_class_meta_field_type_14_is_repeated(q_io_deq_bits_class_meta_field_type_14_is_repeated),
    .io_deq_bits_class_meta_field_type_14_field_type(q_io_deq_bits_class_meta_field_type_14_field_type),
    .io_deq_bits_class_meta_field_type_14_sub_class_id(q_io_deq_bits_class_meta_field_type_14_sub_class_id),
    .io_deq_bits_class_meta_field_type_15_is_repeated(q_io_deq_bits_class_meta_field_type_15_is_repeated),
    .io_deq_bits_class_meta_field_type_15_field_type(q_io_deq_bits_class_meta_field_type_15_field_type),
    .io_deq_bits_class_meta_field_type_15_sub_class_id(q_io_deq_bits_class_meta_field_type_15_sub_class_id),
    .io_deq_bits_class_meta_field_type_16_is_repeated(q_io_deq_bits_class_meta_field_type_16_is_repeated),
    .io_deq_bits_class_meta_field_type_16_field_type(q_io_deq_bits_class_meta_field_type_16_field_type),
    .io_deq_bits_class_meta_field_type_16_sub_class_id(q_io_deq_bits_class_meta_field_type_16_sub_class_id),
    .io_deq_bits_class_meta_field_type_17_is_repeated(q_io_deq_bits_class_meta_field_type_17_is_repeated),
    .io_deq_bits_class_meta_field_type_17_field_type(q_io_deq_bits_class_meta_field_type_17_field_type),
    .io_deq_bits_class_meta_field_type_17_sub_class_id(q_io_deq_bits_class_meta_field_type_17_sub_class_id),
    .io_deq_bits_class_meta_field_type_18_is_repeated(q_io_deq_bits_class_meta_field_type_18_is_repeated),
    .io_deq_bits_class_meta_field_type_18_field_type(q_io_deq_bits_class_meta_field_type_18_field_type),
    .io_deq_bits_class_meta_field_type_18_sub_class_id(q_io_deq_bits_class_meta_field_type_18_sub_class_id),
    .io_deq_bits_class_meta_field_type_19_is_repeated(q_io_deq_bits_class_meta_field_type_19_is_repeated),
    .io_deq_bits_class_meta_field_type_19_field_type(q_io_deq_bits_class_meta_field_type_19_field_type),
    .io_deq_bits_class_meta_field_type_19_sub_class_id(q_io_deq_bits_class_meta_field_type_19_sub_class_id),
    .io_deq_bits_class_meta_field_type_20_is_repeated(q_io_deq_bits_class_meta_field_type_20_is_repeated),
    .io_deq_bits_class_meta_field_type_20_field_type(q_io_deq_bits_class_meta_field_type_20_field_type),
    .io_deq_bits_class_meta_field_type_20_sub_class_id(q_io_deq_bits_class_meta_field_type_20_sub_class_id),
    .io_deq_bits_class_meta_field_type_21_is_repeated(q_io_deq_bits_class_meta_field_type_21_is_repeated),
    .io_deq_bits_class_meta_field_type_21_field_type(q_io_deq_bits_class_meta_field_type_21_field_type),
    .io_deq_bits_class_meta_field_type_21_sub_class_id(q_io_deq_bits_class_meta_field_type_21_sub_class_id),
    .io_deq_bits_class_meta_field_type_22_is_repeated(q_io_deq_bits_class_meta_field_type_22_is_repeated),
    .io_deq_bits_class_meta_field_type_22_field_type(q_io_deq_bits_class_meta_field_type_22_field_type),
    .io_deq_bits_class_meta_field_type_22_sub_class_id(q_io_deq_bits_class_meta_field_type_22_sub_class_id),
    .io_deq_bits_class_meta_field_type_23_is_repeated(q_io_deq_bits_class_meta_field_type_23_is_repeated),
    .io_deq_bits_class_meta_field_type_23_field_type(q_io_deq_bits_class_meta_field_type_23_field_type),
    .io_deq_bits_class_meta_field_type_23_sub_class_id(q_io_deq_bits_class_meta_field_type_23_sub_class_id),
    .io_deq_bits_class_meta_field_type_24_is_repeated(q_io_deq_bits_class_meta_field_type_24_is_repeated),
    .io_deq_bits_class_meta_field_type_24_field_type(q_io_deq_bits_class_meta_field_type_24_field_type),
    .io_deq_bits_class_meta_field_type_24_sub_class_id(q_io_deq_bits_class_meta_field_type_24_sub_class_id),
    .io_deq_bits_class_meta_field_type_25_is_repeated(q_io_deq_bits_class_meta_field_type_25_is_repeated),
    .io_deq_bits_class_meta_field_type_25_field_type(q_io_deq_bits_class_meta_field_type_25_field_type),
    .io_deq_bits_class_meta_field_type_25_sub_class_id(q_io_deq_bits_class_meta_field_type_25_sub_class_id),
    .io_deq_bits_class_meta_field_type_26_is_repeated(q_io_deq_bits_class_meta_field_type_26_is_repeated),
    .io_deq_bits_class_meta_field_type_26_field_type(q_io_deq_bits_class_meta_field_type_26_field_type),
    .io_deq_bits_class_meta_field_type_26_sub_class_id(q_io_deq_bits_class_meta_field_type_26_sub_class_id),
    .io_deq_bits_class_meta_field_type_27_is_repeated(q_io_deq_bits_class_meta_field_type_27_is_repeated),
    .io_deq_bits_class_meta_field_type_27_field_type(q_io_deq_bits_class_meta_field_type_27_field_type),
    .io_deq_bits_class_meta_field_type_27_sub_class_id(q_io_deq_bits_class_meta_field_type_27_sub_class_id),
    .io_deq_bits_class_meta_field_type_28_is_repeated(q_io_deq_bits_class_meta_field_type_28_is_repeated),
    .io_deq_bits_class_meta_field_type_28_field_type(q_io_deq_bits_class_meta_field_type_28_field_type),
    .io_deq_bits_class_meta_field_type_28_sub_class_id(q_io_deq_bits_class_meta_field_type_28_sub_class_id),
    .io_deq_bits_class_meta_field_type_29_is_repeated(q_io_deq_bits_class_meta_field_type_29_is_repeated),
    .io_deq_bits_class_meta_field_type_29_field_type(q_io_deq_bits_class_meta_field_type_29_field_type),
    .io_deq_bits_class_meta_field_type_29_sub_class_id(q_io_deq_bits_class_meta_field_type_29_sub_class_id),
    .io_deq_bits_class_meta_field_type_30_is_repeated(q_io_deq_bits_class_meta_field_type_30_is_repeated),
    .io_deq_bits_class_meta_field_type_30_field_type(q_io_deq_bits_class_meta_field_type_30_field_type),
    .io_deq_bits_class_meta_field_type_30_sub_class_id(q_io_deq_bits_class_meta_field_type_30_sub_class_id),
    .io_deq_bits_class_meta_field_type_31_is_repeated(q_io_deq_bits_class_meta_field_type_31_is_repeated),
    .io_deq_bits_class_meta_field_type_31_field_type(q_io_deq_bits_class_meta_field_type_31_field_type),
    .io_deq_bits_class_meta_field_type_31_sub_class_id(q_io_deq_bits_class_meta_field_type_31_sub_class_id),
    .io_deq_bits_class_meta_field_type_32_is_repeated(q_io_deq_bits_class_meta_field_type_32_is_repeated),
    .io_deq_bits_class_meta_field_type_32_field_type(q_io_deq_bits_class_meta_field_type_32_field_type),
    .io_deq_bits_class_meta_field_type_32_sub_class_id(q_io_deq_bits_class_meta_field_type_32_sub_class_id)
  );
  assign io_out_valid = q_io_deq_valid; // @[XQueue.scala 88:34]
  assign io_out_bits_class_meta_max_field_num = q_io_deq_bits_class_meta_max_field_num; // @[XQueue.scala 88:34]
  assign io_out_bits_class_meta_field_type_0_is_repeated = q_io_deq_bits_class_meta_field_type_0_is_repeated; // @[XQueue.scala 88:34]
  assign io_out_bits_class_meta_field_type_0_field_type = q_io_deq_bits_class_meta_field_type_0_field_type; // @[XQueue.scala 88:34]
  assign io_out_bits_class_meta_field_type_0_sub_class_id = q_io_deq_bits_class_meta_field_type_0_sub_class_id; // @[XQueue.scala 88:34]
  assign io_out_bits_class_meta_field_type_1_is_repeated = q_io_deq_bits_class_meta_field_type_1_is_repeated; // @[XQueue.scala 88:34]
  assign io_out_bits_class_meta_field_type_1_field_type = q_io_deq_bits_class_meta_field_type_1_field_type; // @[XQueue.scala 88:34]
  assign io_out_bits_class_meta_field_type_1_sub_class_id = q_io_deq_bits_class_meta_field_type_1_sub_class_id; // @[XQueue.scala 88:34]
  assign io_out_bits_class_meta_field_type_2_is_repeated = q_io_deq_bits_class_meta_field_type_2_is_repeated; // @[XQueue.scala 88:34]
  assign io_out_bits_class_meta_field_type_2_field_type = q_io_deq_bits_class_meta_field_type_2_field_type; // @[XQueue.scala 88:34]
  assign io_out_bits_class_meta_field_type_2_sub_class_id = q_io_deq_bits_class_meta_field_type_2_sub_class_id; // @[XQueue.scala 88:34]
  assign io_out_bits_class_meta_field_type_3_is_repeated = q_io_deq_bits_class_meta_field_type_3_is_repeated; // @[XQueue.scala 88:34]
  assign io_out_bits_class_meta_field_type_3_field_type = q_io_deq_bits_class_meta_field_type_3_field_type; // @[XQueue.scala 88:34]
  assign io_out_bits_class_meta_field_type_3_sub_class_id = q_io_deq_bits_class_meta_field_type_3_sub_class_id; // @[XQueue.scala 88:34]
  assign io_out_bits_class_meta_field_type_4_is_repeated = q_io_deq_bits_class_meta_field_type_4_is_repeated; // @[XQueue.scala 88:34]
  assign io_out_bits_class_meta_field_type_4_field_type = q_io_deq_bits_class_meta_field_type_4_field_type; // @[XQueue.scala 88:34]
  assign io_out_bits_class_meta_field_type_4_sub_class_id = q_io_deq_bits_class_meta_field_type_4_sub_class_id; // @[XQueue.scala 88:34]
  assign io_out_bits_class_meta_field_type_5_is_repeated = q_io_deq_bits_class_meta_field_type_5_is_repeated; // @[XQueue.scala 88:34]
  assign io_out_bits_class_meta_field_type_5_field_type = q_io_deq_bits_class_meta_field_type_5_field_type; // @[XQueue.scala 88:34]
  assign io_out_bits_class_meta_field_type_5_sub_class_id = q_io_deq_bits_class_meta_field_type_5_sub_class_id; // @[XQueue.scala 88:34]
  assign io_out_bits_class_meta_field_type_6_is_repeated = q_io_deq_bits_class_meta_field_type_6_is_repeated; // @[XQueue.scala 88:34]
  assign io_out_bits_class_meta_field_type_6_field_type = q_io_deq_bits_class_meta_field_type_6_field_type; // @[XQueue.scala 88:34]
  assign io_out_bits_class_meta_field_type_6_sub_class_id = q_io_deq_bits_class_meta_field_type_6_sub_class_id; // @[XQueue.scala 88:34]
  assign io_out_bits_class_meta_field_type_7_is_repeated = q_io_deq_bits_class_meta_field_type_7_is_repeated; // @[XQueue.scala 88:34]
  assign io_out_bits_class_meta_field_type_7_field_type = q_io_deq_bits_class_meta_field_type_7_field_type; // @[XQueue.scala 88:34]
  assign io_out_bits_class_meta_field_type_7_sub_class_id = q_io_deq_bits_class_meta_field_type_7_sub_class_id; // @[XQueue.scala 88:34]
  assign io_out_bits_class_meta_field_type_8_is_repeated = q_io_deq_bits_class_meta_field_type_8_is_repeated; // @[XQueue.scala 88:34]
  assign io_out_bits_class_meta_field_type_8_field_type = q_io_deq_bits_class_meta_field_type_8_field_type; // @[XQueue.scala 88:34]
  assign io_out_bits_class_meta_field_type_8_sub_class_id = q_io_deq_bits_class_meta_field_type_8_sub_class_id; // @[XQueue.scala 88:34]
  assign io_out_bits_class_meta_field_type_9_is_repeated = q_io_deq_bits_class_meta_field_type_9_is_repeated; // @[XQueue.scala 88:34]
  assign io_out_bits_class_meta_field_type_9_field_type = q_io_deq_bits_class_meta_field_type_9_field_type; // @[XQueue.scala 88:34]
  assign io_out_bits_class_meta_field_type_9_sub_class_id = q_io_deq_bits_class_meta_field_type_9_sub_class_id; // @[XQueue.scala 88:34]
  assign io_out_bits_class_meta_field_type_10_is_repeated = q_io_deq_bits_class_meta_field_type_10_is_repeated; // @[XQueue.scala 88:34]
  assign io_out_bits_class_meta_field_type_10_field_type = q_io_deq_bits_class_meta_field_type_10_field_type; // @[XQueue.scala 88:34]
  assign io_out_bits_class_meta_field_type_10_sub_class_id = q_io_deq_bits_class_meta_field_type_10_sub_class_id; // @[XQueue.scala 88:34]
  assign io_out_bits_class_meta_field_type_11_is_repeated = q_io_deq_bits_class_meta_field_type_11_is_repeated; // @[XQueue.scala 88:34]
  assign io_out_bits_class_meta_field_type_11_field_type = q_io_deq_bits_class_meta_field_type_11_field_type; // @[XQueue.scala 88:34]
  assign io_out_bits_class_meta_field_type_11_sub_class_id = q_io_deq_bits_class_meta_field_type_11_sub_class_id; // @[XQueue.scala 88:34]
  assign io_out_bits_class_meta_field_type_12_is_repeated = q_io_deq_bits_class_meta_field_type_12_is_repeated; // @[XQueue.scala 88:34]
  assign io_out_bits_class_meta_field_type_12_field_type = q_io_deq_bits_class_meta_field_type_12_field_type; // @[XQueue.scala 88:34]
  assign io_out_bits_class_meta_field_type_12_sub_class_id = q_io_deq_bits_class_meta_field_type_12_sub_class_id; // @[XQueue.scala 88:34]
  assign io_out_bits_class_meta_field_type_13_is_repeated = q_io_deq_bits_class_meta_field_type_13_is_repeated; // @[XQueue.scala 88:34]
  assign io_out_bits_class_meta_field_type_13_field_type = q_io_deq_bits_class_meta_field_type_13_field_type; // @[XQueue.scala 88:34]
  assign io_out_bits_class_meta_field_type_13_sub_class_id = q_io_deq_bits_class_meta_field_type_13_sub_class_id; // @[XQueue.scala 88:34]
  assign io_out_bits_class_meta_field_type_14_is_repeated = q_io_deq_bits_class_meta_field_type_14_is_repeated; // @[XQueue.scala 88:34]
  assign io_out_bits_class_meta_field_type_14_field_type = q_io_deq_bits_class_meta_field_type_14_field_type; // @[XQueue.scala 88:34]
  assign io_out_bits_class_meta_field_type_14_sub_class_id = q_io_deq_bits_class_meta_field_type_14_sub_class_id; // @[XQueue.scala 88:34]
  assign io_out_bits_class_meta_field_type_15_is_repeated = q_io_deq_bits_class_meta_field_type_15_is_repeated; // @[XQueue.scala 88:34]
  assign io_out_bits_class_meta_field_type_15_field_type = q_io_deq_bits_class_meta_field_type_15_field_type; // @[XQueue.scala 88:34]
  assign io_out_bits_class_meta_field_type_15_sub_class_id = q_io_deq_bits_class_meta_field_type_15_sub_class_id; // @[XQueue.scala 88:34]
  assign io_out_bits_class_meta_field_type_16_is_repeated = q_io_deq_bits_class_meta_field_type_16_is_repeated; // @[XQueue.scala 88:34]
  assign io_out_bits_class_meta_field_type_16_field_type = q_io_deq_bits_class_meta_field_type_16_field_type; // @[XQueue.scala 88:34]
  assign io_out_bits_class_meta_field_type_16_sub_class_id = q_io_deq_bits_class_meta_field_type_16_sub_class_id; // @[XQueue.scala 88:34]
  assign io_out_bits_class_meta_field_type_17_is_repeated = q_io_deq_bits_class_meta_field_type_17_is_repeated; // @[XQueue.scala 88:34]
  assign io_out_bits_class_meta_field_type_17_field_type = q_io_deq_bits_class_meta_field_type_17_field_type; // @[XQueue.scala 88:34]
  assign io_out_bits_class_meta_field_type_17_sub_class_id = q_io_deq_bits_class_meta_field_type_17_sub_class_id; // @[XQueue.scala 88:34]
  assign io_out_bits_class_meta_field_type_18_is_repeated = q_io_deq_bits_class_meta_field_type_18_is_repeated; // @[XQueue.scala 88:34]
  assign io_out_bits_class_meta_field_type_18_field_type = q_io_deq_bits_class_meta_field_type_18_field_type; // @[XQueue.scala 88:34]
  assign io_out_bits_class_meta_field_type_18_sub_class_id = q_io_deq_bits_class_meta_field_type_18_sub_class_id; // @[XQueue.scala 88:34]
  assign io_out_bits_class_meta_field_type_19_is_repeated = q_io_deq_bits_class_meta_field_type_19_is_repeated; // @[XQueue.scala 88:34]
  assign io_out_bits_class_meta_field_type_19_field_type = q_io_deq_bits_class_meta_field_type_19_field_type; // @[XQueue.scala 88:34]
  assign io_out_bits_class_meta_field_type_19_sub_class_id = q_io_deq_bits_class_meta_field_type_19_sub_class_id; // @[XQueue.scala 88:34]
  assign io_out_bits_class_meta_field_type_20_is_repeated = q_io_deq_bits_class_meta_field_type_20_is_repeated; // @[XQueue.scala 88:34]
  assign io_out_bits_class_meta_field_type_20_field_type = q_io_deq_bits_class_meta_field_type_20_field_type; // @[XQueue.scala 88:34]
  assign io_out_bits_class_meta_field_type_20_sub_class_id = q_io_deq_bits_class_meta_field_type_20_sub_class_id; // @[XQueue.scala 88:34]
  assign io_out_bits_class_meta_field_type_21_is_repeated = q_io_deq_bits_class_meta_field_type_21_is_repeated; // @[XQueue.scala 88:34]
  assign io_out_bits_class_meta_field_type_21_field_type = q_io_deq_bits_class_meta_field_type_21_field_type; // @[XQueue.scala 88:34]
  assign io_out_bits_class_meta_field_type_21_sub_class_id = q_io_deq_bits_class_meta_field_type_21_sub_class_id; // @[XQueue.scala 88:34]
  assign io_out_bits_class_meta_field_type_22_is_repeated = q_io_deq_bits_class_meta_field_type_22_is_repeated; // @[XQueue.scala 88:34]
  assign io_out_bits_class_meta_field_type_22_field_type = q_io_deq_bits_class_meta_field_type_22_field_type; // @[XQueue.scala 88:34]
  assign io_out_bits_class_meta_field_type_22_sub_class_id = q_io_deq_bits_class_meta_field_type_22_sub_class_id; // @[XQueue.scala 88:34]
  assign io_out_bits_class_meta_field_type_23_is_repeated = q_io_deq_bits_class_meta_field_type_23_is_repeated; // @[XQueue.scala 88:34]
  assign io_out_bits_class_meta_field_type_23_field_type = q_io_deq_bits_class_meta_field_type_23_field_type; // @[XQueue.scala 88:34]
  assign io_out_bits_class_meta_field_type_23_sub_class_id = q_io_deq_bits_class_meta_field_type_23_sub_class_id; // @[XQueue.scala 88:34]
  assign io_out_bits_class_meta_field_type_24_is_repeated = q_io_deq_bits_class_meta_field_type_24_is_repeated; // @[XQueue.scala 88:34]
  assign io_out_bits_class_meta_field_type_24_field_type = q_io_deq_bits_class_meta_field_type_24_field_type; // @[XQueue.scala 88:34]
  assign io_out_bits_class_meta_field_type_24_sub_class_id = q_io_deq_bits_class_meta_field_type_24_sub_class_id; // @[XQueue.scala 88:34]
  assign io_out_bits_class_meta_field_type_25_is_repeated = q_io_deq_bits_class_meta_field_type_25_is_repeated; // @[XQueue.scala 88:34]
  assign io_out_bits_class_meta_field_type_25_field_type = q_io_deq_bits_class_meta_field_type_25_field_type; // @[XQueue.scala 88:34]
  assign io_out_bits_class_meta_field_type_25_sub_class_id = q_io_deq_bits_class_meta_field_type_25_sub_class_id; // @[XQueue.scala 88:34]
  assign io_out_bits_class_meta_field_type_26_is_repeated = q_io_deq_bits_class_meta_field_type_26_is_repeated; // @[XQueue.scala 88:34]
  assign io_out_bits_class_meta_field_type_26_field_type = q_io_deq_bits_class_meta_field_type_26_field_type; // @[XQueue.scala 88:34]
  assign io_out_bits_class_meta_field_type_26_sub_class_id = q_io_deq_bits_class_meta_field_type_26_sub_class_id; // @[XQueue.scala 88:34]
  assign io_out_bits_class_meta_field_type_27_is_repeated = q_io_deq_bits_class_meta_field_type_27_is_repeated; // @[XQueue.scala 88:34]
  assign io_out_bits_class_meta_field_type_27_field_type = q_io_deq_bits_class_meta_field_type_27_field_type; // @[XQueue.scala 88:34]
  assign io_out_bits_class_meta_field_type_27_sub_class_id = q_io_deq_bits_class_meta_field_type_27_sub_class_id; // @[XQueue.scala 88:34]
  assign io_out_bits_class_meta_field_type_28_is_repeated = q_io_deq_bits_class_meta_field_type_28_is_repeated; // @[XQueue.scala 88:34]
  assign io_out_bits_class_meta_field_type_28_field_type = q_io_deq_bits_class_meta_field_type_28_field_type; // @[XQueue.scala 88:34]
  assign io_out_bits_class_meta_field_type_28_sub_class_id = q_io_deq_bits_class_meta_field_type_28_sub_class_id; // @[XQueue.scala 88:34]
  assign io_out_bits_class_meta_field_type_29_is_repeated = q_io_deq_bits_class_meta_field_type_29_is_repeated; // @[XQueue.scala 88:34]
  assign io_out_bits_class_meta_field_type_29_field_type = q_io_deq_bits_class_meta_field_type_29_field_type; // @[XQueue.scala 88:34]
  assign io_out_bits_class_meta_field_type_29_sub_class_id = q_io_deq_bits_class_meta_field_type_29_sub_class_id; // @[XQueue.scala 88:34]
  assign io_out_bits_class_meta_field_type_30_is_repeated = q_io_deq_bits_class_meta_field_type_30_is_repeated; // @[XQueue.scala 88:34]
  assign io_out_bits_class_meta_field_type_30_field_type = q_io_deq_bits_class_meta_field_type_30_field_type; // @[XQueue.scala 88:34]
  assign io_out_bits_class_meta_field_type_30_sub_class_id = q_io_deq_bits_class_meta_field_type_30_sub_class_id; // @[XQueue.scala 88:34]
  assign io_out_bits_class_meta_field_type_31_is_repeated = q_io_deq_bits_class_meta_field_type_31_is_repeated; // @[XQueue.scala 88:34]
  assign io_out_bits_class_meta_field_type_31_field_type = q_io_deq_bits_class_meta_field_type_31_field_type; // @[XQueue.scala 88:34]
  assign io_out_bits_class_meta_field_type_31_sub_class_id = q_io_deq_bits_class_meta_field_type_31_sub_class_id; // @[XQueue.scala 88:34]
  assign io_out_bits_class_meta_field_type_32_is_repeated = q_io_deq_bits_class_meta_field_type_32_is_repeated; // @[XQueue.scala 88:34]
  assign io_out_bits_class_meta_field_type_32_field_type = q_io_deq_bits_class_meta_field_type_32_field_type; // @[XQueue.scala 88:34]
  assign io_out_bits_class_meta_field_type_32_sub_class_id = q_io_deq_bits_class_meta_field_type_32_sub_class_id; // @[XQueue.scala 88:34]
  assign q_clock = clock;
  assign q_reset = reset;
  assign q_io_enq_valid = io_in_valid; // @[XQueue.scala 87:34]
  assign q_io_enq_bits_class_meta_max_field_num = io_in_bits_class_meta_max_field_num; // @[XQueue.scala 87:34]
  assign q_io_enq_bits_class_meta_field_type_0_is_repeated = io_in_bits_class_meta_field_type_0_is_repeated; // @[XQueue.scala 87:34]
  assign q_io_enq_bits_class_meta_field_type_0_field_type = io_in_bits_class_meta_field_type_0_field_type; // @[XQueue.scala 87:34]
  assign q_io_enq_bits_class_meta_field_type_0_sub_class_id = io_in_bits_class_meta_field_type_0_sub_class_id; // @[XQueue.scala 87:34]
  assign q_io_enq_bits_class_meta_field_type_1_is_repeated = io_in_bits_class_meta_field_type_1_is_repeated; // @[XQueue.scala 87:34]
  assign q_io_enq_bits_class_meta_field_type_1_field_type = io_in_bits_class_meta_field_type_1_field_type; // @[XQueue.scala 87:34]
  assign q_io_enq_bits_class_meta_field_type_1_sub_class_id = io_in_bits_class_meta_field_type_1_sub_class_id; // @[XQueue.scala 87:34]
  assign q_io_enq_bits_class_meta_field_type_2_is_repeated = io_in_bits_class_meta_field_type_2_is_repeated; // @[XQueue.scala 87:34]
  assign q_io_enq_bits_class_meta_field_type_2_field_type = io_in_bits_class_meta_field_type_2_field_type; // @[XQueue.scala 87:34]
  assign q_io_enq_bits_class_meta_field_type_2_sub_class_id = io_in_bits_class_meta_field_type_2_sub_class_id; // @[XQueue.scala 87:34]
  assign q_io_enq_bits_class_meta_field_type_3_is_repeated = io_in_bits_class_meta_field_type_3_is_repeated; // @[XQueue.scala 87:34]
  assign q_io_enq_bits_class_meta_field_type_3_field_type = io_in_bits_class_meta_field_type_3_field_type; // @[XQueue.scala 87:34]
  assign q_io_enq_bits_class_meta_field_type_3_sub_class_id = io_in_bits_class_meta_field_type_3_sub_class_id; // @[XQueue.scala 87:34]
  assign q_io_enq_bits_class_meta_field_type_4_is_repeated = io_in_bits_class_meta_field_type_4_is_repeated; // @[XQueue.scala 87:34]
  assign q_io_enq_bits_class_meta_field_type_4_field_type = io_in_bits_class_meta_field_type_4_field_type; // @[XQueue.scala 87:34]
  assign q_io_enq_bits_class_meta_field_type_4_sub_class_id = io_in_bits_class_meta_field_type_4_sub_class_id; // @[XQueue.scala 87:34]
  assign q_io_enq_bits_class_meta_field_type_5_is_repeated = io_in_bits_class_meta_field_type_5_is_repeated; // @[XQueue.scala 87:34]
  assign q_io_enq_bits_class_meta_field_type_5_field_type = io_in_bits_class_meta_field_type_5_field_type; // @[XQueue.scala 87:34]
  assign q_io_enq_bits_class_meta_field_type_5_sub_class_id = io_in_bits_class_meta_field_type_5_sub_class_id; // @[XQueue.scala 87:34]
  assign q_io_enq_bits_class_meta_field_type_6_is_repeated = io_in_bits_class_meta_field_type_6_is_repeated; // @[XQueue.scala 87:34]
  assign q_io_enq_bits_class_meta_field_type_6_field_type = io_in_bits_class_meta_field_type_6_field_type; // @[XQueue.scala 87:34]
  assign q_io_enq_bits_class_meta_field_type_6_sub_class_id = io_in_bits_class_meta_field_type_6_sub_class_id; // @[XQueue.scala 87:34]
  assign q_io_enq_bits_class_meta_field_type_7_is_repeated = io_in_bits_class_meta_field_type_7_is_repeated; // @[XQueue.scala 87:34]
  assign q_io_enq_bits_class_meta_field_type_7_field_type = io_in_bits_class_meta_field_type_7_field_type; // @[XQueue.scala 87:34]
  assign q_io_enq_bits_class_meta_field_type_7_sub_class_id = io_in_bits_class_meta_field_type_7_sub_class_id; // @[XQueue.scala 87:34]
  assign q_io_enq_bits_class_meta_field_type_8_is_repeated = io_in_bits_class_meta_field_type_8_is_repeated; // @[XQueue.scala 87:34]
  assign q_io_enq_bits_class_meta_field_type_8_field_type = io_in_bits_class_meta_field_type_8_field_type; // @[XQueue.scala 87:34]
  assign q_io_enq_bits_class_meta_field_type_8_sub_class_id = io_in_bits_class_meta_field_type_8_sub_class_id; // @[XQueue.scala 87:34]
  assign q_io_enq_bits_class_meta_field_type_9_is_repeated = io_in_bits_class_meta_field_type_9_is_repeated; // @[XQueue.scala 87:34]
  assign q_io_enq_bits_class_meta_field_type_9_field_type = io_in_bits_class_meta_field_type_9_field_type; // @[XQueue.scala 87:34]
  assign q_io_enq_bits_class_meta_field_type_9_sub_class_id = io_in_bits_class_meta_field_type_9_sub_class_id; // @[XQueue.scala 87:34]
  assign q_io_enq_bits_class_meta_field_type_10_is_repeated = io_in_bits_class_meta_field_type_10_is_repeated; // @[XQueue.scala 87:34]
  assign q_io_enq_bits_class_meta_field_type_10_field_type = io_in_bits_class_meta_field_type_10_field_type; // @[XQueue.scala 87:34]
  assign q_io_enq_bits_class_meta_field_type_10_sub_class_id = io_in_bits_class_meta_field_type_10_sub_class_id; // @[XQueue.scala 87:34]
  assign q_io_enq_bits_class_meta_field_type_11_is_repeated = io_in_bits_class_meta_field_type_11_is_repeated; // @[XQueue.scala 87:34]
  assign q_io_enq_bits_class_meta_field_type_11_field_type = io_in_bits_class_meta_field_type_11_field_type; // @[XQueue.scala 87:34]
  assign q_io_enq_bits_class_meta_field_type_11_sub_class_id = io_in_bits_class_meta_field_type_11_sub_class_id; // @[XQueue.scala 87:34]
  assign q_io_enq_bits_class_meta_field_type_12_is_repeated = io_in_bits_class_meta_field_type_12_is_repeated; // @[XQueue.scala 87:34]
  assign q_io_enq_bits_class_meta_field_type_12_field_type = io_in_bits_class_meta_field_type_12_field_type; // @[XQueue.scala 87:34]
  assign q_io_enq_bits_class_meta_field_type_12_sub_class_id = io_in_bits_class_meta_field_type_12_sub_class_id; // @[XQueue.scala 87:34]
  assign q_io_enq_bits_class_meta_field_type_13_is_repeated = io_in_bits_class_meta_field_type_13_is_repeated; // @[XQueue.scala 87:34]
  assign q_io_enq_bits_class_meta_field_type_13_field_type = io_in_bits_class_meta_field_type_13_field_type; // @[XQueue.scala 87:34]
  assign q_io_enq_bits_class_meta_field_type_13_sub_class_id = io_in_bits_class_meta_field_type_13_sub_class_id; // @[XQueue.scala 87:34]
  assign q_io_enq_bits_class_meta_field_type_14_is_repeated = io_in_bits_class_meta_field_type_14_is_repeated; // @[XQueue.scala 87:34]
  assign q_io_enq_bits_class_meta_field_type_14_field_type = io_in_bits_class_meta_field_type_14_field_type; // @[XQueue.scala 87:34]
  assign q_io_enq_bits_class_meta_field_type_14_sub_class_id = io_in_bits_class_meta_field_type_14_sub_class_id; // @[XQueue.scala 87:34]
  assign q_io_enq_bits_class_meta_field_type_15_is_repeated = io_in_bits_class_meta_field_type_15_is_repeated; // @[XQueue.scala 87:34]
  assign q_io_enq_bits_class_meta_field_type_15_field_type = io_in_bits_class_meta_field_type_15_field_type; // @[XQueue.scala 87:34]
  assign q_io_enq_bits_class_meta_field_type_15_sub_class_id = io_in_bits_class_meta_field_type_15_sub_class_id; // @[XQueue.scala 87:34]
  assign q_io_enq_bits_class_meta_field_type_16_is_repeated = io_in_bits_class_meta_field_type_16_is_repeated; // @[XQueue.scala 87:34]
  assign q_io_enq_bits_class_meta_field_type_16_field_type = io_in_bits_class_meta_field_type_16_field_type; // @[XQueue.scala 87:34]
  assign q_io_enq_bits_class_meta_field_type_16_sub_class_id = io_in_bits_class_meta_field_type_16_sub_class_id; // @[XQueue.scala 87:34]
  assign q_io_enq_bits_class_meta_field_type_17_is_repeated = io_in_bits_class_meta_field_type_17_is_repeated; // @[XQueue.scala 87:34]
  assign q_io_enq_bits_class_meta_field_type_17_field_type = io_in_bits_class_meta_field_type_17_field_type; // @[XQueue.scala 87:34]
  assign q_io_enq_bits_class_meta_field_type_17_sub_class_id = io_in_bits_class_meta_field_type_17_sub_class_id; // @[XQueue.scala 87:34]
  assign q_io_enq_bits_class_meta_field_type_18_is_repeated = io_in_bits_class_meta_field_type_18_is_repeated; // @[XQueue.scala 87:34]
  assign q_io_enq_bits_class_meta_field_type_18_field_type = io_in_bits_class_meta_field_type_18_field_type; // @[XQueue.scala 87:34]
  assign q_io_enq_bits_class_meta_field_type_18_sub_class_id = io_in_bits_class_meta_field_type_18_sub_class_id; // @[XQueue.scala 87:34]
  assign q_io_enq_bits_class_meta_field_type_19_is_repeated = io_in_bits_class_meta_field_type_19_is_repeated; // @[XQueue.scala 87:34]
  assign q_io_enq_bits_class_meta_field_type_19_field_type = io_in_bits_class_meta_field_type_19_field_type; // @[XQueue.scala 87:34]
  assign q_io_enq_bits_class_meta_field_type_19_sub_class_id = io_in_bits_class_meta_field_type_19_sub_class_id; // @[XQueue.scala 87:34]
  assign q_io_enq_bits_class_meta_field_type_20_is_repeated = io_in_bits_class_meta_field_type_20_is_repeated; // @[XQueue.scala 87:34]
  assign q_io_enq_bits_class_meta_field_type_20_field_type = io_in_bits_class_meta_field_type_20_field_type; // @[XQueue.scala 87:34]
  assign q_io_enq_bits_class_meta_field_type_20_sub_class_id = io_in_bits_class_meta_field_type_20_sub_class_id; // @[XQueue.scala 87:34]
  assign q_io_enq_bits_class_meta_field_type_21_is_repeated = io_in_bits_class_meta_field_type_21_is_repeated; // @[XQueue.scala 87:34]
  assign q_io_enq_bits_class_meta_field_type_21_field_type = io_in_bits_class_meta_field_type_21_field_type; // @[XQueue.scala 87:34]
  assign q_io_enq_bits_class_meta_field_type_21_sub_class_id = io_in_bits_class_meta_field_type_21_sub_class_id; // @[XQueue.scala 87:34]
  assign q_io_enq_bits_class_meta_field_type_22_is_repeated = io_in_bits_class_meta_field_type_22_is_repeated; // @[XQueue.scala 87:34]
  assign q_io_enq_bits_class_meta_field_type_22_field_type = io_in_bits_class_meta_field_type_22_field_type; // @[XQueue.scala 87:34]
  assign q_io_enq_bits_class_meta_field_type_22_sub_class_id = io_in_bits_class_meta_field_type_22_sub_class_id; // @[XQueue.scala 87:34]
  assign q_io_enq_bits_class_meta_field_type_23_is_repeated = io_in_bits_class_meta_field_type_23_is_repeated; // @[XQueue.scala 87:34]
  assign q_io_enq_bits_class_meta_field_type_23_field_type = io_in_bits_class_meta_field_type_23_field_type; // @[XQueue.scala 87:34]
  assign q_io_enq_bits_class_meta_field_type_23_sub_class_id = io_in_bits_class_meta_field_type_23_sub_class_id; // @[XQueue.scala 87:34]
  assign q_io_enq_bits_class_meta_field_type_24_is_repeated = io_in_bits_class_meta_field_type_24_is_repeated; // @[XQueue.scala 87:34]
  assign q_io_enq_bits_class_meta_field_type_24_field_type = io_in_bits_class_meta_field_type_24_field_type; // @[XQueue.scala 87:34]
  assign q_io_enq_bits_class_meta_field_type_24_sub_class_id = io_in_bits_class_meta_field_type_24_sub_class_id; // @[XQueue.scala 87:34]
  assign q_io_enq_bits_class_meta_field_type_25_is_repeated = io_in_bits_class_meta_field_type_25_is_repeated; // @[XQueue.scala 87:34]
  assign q_io_enq_bits_class_meta_field_type_25_field_type = io_in_bits_class_meta_field_type_25_field_type; // @[XQueue.scala 87:34]
  assign q_io_enq_bits_class_meta_field_type_25_sub_class_id = io_in_bits_class_meta_field_type_25_sub_class_id; // @[XQueue.scala 87:34]
  assign q_io_enq_bits_class_meta_field_type_26_is_repeated = io_in_bits_class_meta_field_type_26_is_repeated; // @[XQueue.scala 87:34]
  assign q_io_enq_bits_class_meta_field_type_26_field_type = io_in_bits_class_meta_field_type_26_field_type; // @[XQueue.scala 87:34]
  assign q_io_enq_bits_class_meta_field_type_26_sub_class_id = io_in_bits_class_meta_field_type_26_sub_class_id; // @[XQueue.scala 87:34]
  assign q_io_enq_bits_class_meta_field_type_27_is_repeated = io_in_bits_class_meta_field_type_27_is_repeated; // @[XQueue.scala 87:34]
  assign q_io_enq_bits_class_meta_field_type_27_field_type = io_in_bits_class_meta_field_type_27_field_type; // @[XQueue.scala 87:34]
  assign q_io_enq_bits_class_meta_field_type_27_sub_class_id = io_in_bits_class_meta_field_type_27_sub_class_id; // @[XQueue.scala 87:34]
  assign q_io_enq_bits_class_meta_field_type_28_is_repeated = io_in_bits_class_meta_field_type_28_is_repeated; // @[XQueue.scala 87:34]
  assign q_io_enq_bits_class_meta_field_type_28_field_type = io_in_bits_class_meta_field_type_28_field_type; // @[XQueue.scala 87:34]
  assign q_io_enq_bits_class_meta_field_type_28_sub_class_id = io_in_bits_class_meta_field_type_28_sub_class_id; // @[XQueue.scala 87:34]
  assign q_io_enq_bits_class_meta_field_type_29_is_repeated = io_in_bits_class_meta_field_type_29_is_repeated; // @[XQueue.scala 87:34]
  assign q_io_enq_bits_class_meta_field_type_29_field_type = io_in_bits_class_meta_field_type_29_field_type; // @[XQueue.scala 87:34]
  assign q_io_enq_bits_class_meta_field_type_29_sub_class_id = io_in_bits_class_meta_field_type_29_sub_class_id; // @[XQueue.scala 87:34]
  assign q_io_enq_bits_class_meta_field_type_30_is_repeated = io_in_bits_class_meta_field_type_30_is_repeated; // @[XQueue.scala 87:34]
  assign q_io_enq_bits_class_meta_field_type_30_field_type = io_in_bits_class_meta_field_type_30_field_type; // @[XQueue.scala 87:34]
  assign q_io_enq_bits_class_meta_field_type_30_sub_class_id = io_in_bits_class_meta_field_type_30_sub_class_id; // @[XQueue.scala 87:34]
  assign q_io_enq_bits_class_meta_field_type_31_is_repeated = io_in_bits_class_meta_field_type_31_is_repeated; // @[XQueue.scala 87:34]
  assign q_io_enq_bits_class_meta_field_type_31_field_type = io_in_bits_class_meta_field_type_31_field_type; // @[XQueue.scala 87:34]
  assign q_io_enq_bits_class_meta_field_type_31_sub_class_id = io_in_bits_class_meta_field_type_31_sub_class_id; // @[XQueue.scala 87:34]
  assign q_io_enq_bits_class_meta_field_type_32_is_repeated = io_in_bits_class_meta_field_type_32_is_repeated; // @[XQueue.scala 87:34]
  assign q_io_enq_bits_class_meta_field_type_32_field_type = io_in_bits_class_meta_field_type_32_field_type; // @[XQueue.scala 87:34]
  assign q_io_enq_bits_class_meta_field_type_32_sub_class_id = io_in_bits_class_meta_field_type_32_sub_class_id; // @[XQueue.scala 87:34]
  assign q_io_deq_ready = io_out_ready; // @[XQueue.scala 88:34]
endmodule
module Serializerhw(
  input         clock,
  input         reset,
  output        io_meta_in_ready,
  input         io_meta_in_valid,
  input  [9:0]  io_meta_in_bits_class_id,
  input  [63:0] io_meta_in_bits_host_base_addr,
  output        io_host_data_in_ready,
  input         io_host_data_in_valid,
  input         io_host_data_cmd_ready,
  output        io_host_data_cmd_valid,
  output [63:0] io_host_data_cmd_bits_vaddr,
  output [31:0] io_host_data_cmd_bits_length,
  input         io_class_meta_req_ready,
  output        io_class_meta_req_valid,
  output [9:0]  io_class_meta_req_bits_class_id,
  input         io_class_meta_rsp_valid,
  input  [7:0]  io_class_meta_rsp_bits_class_meta_max_field_num,
  input         io_class_meta_rsp_bits_class_meta_field_type_0_is_repeated,
  input  [4:0]  io_class_meta_rsp_bits_class_meta_field_type_0_field_type,
  input  [15:0] io_class_meta_rsp_bits_class_meta_field_type_0_sub_class_id,
  input         io_class_meta_rsp_bits_class_meta_field_type_1_is_repeated,
  input  [4:0]  io_class_meta_rsp_bits_class_meta_field_type_1_field_type,
  input  [15:0] io_class_meta_rsp_bits_class_meta_field_type_1_sub_class_id,
  input         io_class_meta_rsp_bits_class_meta_field_type_2_is_repeated,
  input  [4:0]  io_class_meta_rsp_bits_class_meta_field_type_2_field_type,
  input  [15:0] io_class_meta_rsp_bits_class_meta_field_type_2_sub_class_id,
  input         io_class_meta_rsp_bits_class_meta_field_type_3_is_repeated,
  input  [4:0]  io_class_meta_rsp_bits_class_meta_field_type_3_field_type,
  input  [15:0] io_class_meta_rsp_bits_class_meta_field_type_3_sub_class_id,
  input         io_class_meta_rsp_bits_class_meta_field_type_4_is_repeated,
  input  [4:0]  io_class_meta_rsp_bits_class_meta_field_type_4_field_type,
  input  [15:0] io_class_meta_rsp_bits_class_meta_field_type_4_sub_class_id,
  input         io_class_meta_rsp_bits_class_meta_field_type_5_is_repeated,
  input  [4:0]  io_class_meta_rsp_bits_class_meta_field_type_5_field_type,
  input  [15:0] io_class_meta_rsp_bits_class_meta_field_type_5_sub_class_id,
  input         io_class_meta_rsp_bits_class_meta_field_type_6_is_repeated,
  input  [4:0]  io_class_meta_rsp_bits_class_meta_field_type_6_field_type,
  input  [15:0] io_class_meta_rsp_bits_class_meta_field_type_6_sub_class_id,
  input         io_class_meta_rsp_bits_class_meta_field_type_7_is_repeated,
  input  [4:0]  io_class_meta_rsp_bits_class_meta_field_type_7_field_type,
  input  [15:0] io_class_meta_rsp_bits_class_meta_field_type_7_sub_class_id,
  input         io_class_meta_rsp_bits_class_meta_field_type_8_is_repeated,
  input  [4:0]  io_class_meta_rsp_bits_class_meta_field_type_8_field_type,
  input  [15:0] io_class_meta_rsp_bits_class_meta_field_type_8_sub_class_id,
  input         io_class_meta_rsp_bits_class_meta_field_type_9_is_repeated,
  input  [4:0]  io_class_meta_rsp_bits_class_meta_field_type_9_field_type,
  input  [15:0] io_class_meta_rsp_bits_class_meta_field_type_9_sub_class_id,
  input         io_class_meta_rsp_bits_class_meta_field_type_10_is_repeated,
  input  [4:0]  io_class_meta_rsp_bits_class_meta_field_type_10_field_type,
  input  [15:0] io_class_meta_rsp_bits_class_meta_field_type_10_sub_class_id,
  input         io_class_meta_rsp_bits_class_meta_field_type_11_is_repeated,
  input  [4:0]  io_class_meta_rsp_bits_class_meta_field_type_11_field_type,
  input  [15:0] io_class_meta_rsp_bits_class_meta_field_type_11_sub_class_id,
  input         io_class_meta_rsp_bits_class_meta_field_type_12_is_repeated,
  input  [4:0]  io_class_meta_rsp_bits_class_meta_field_type_12_field_type,
  input  [15:0] io_class_meta_rsp_bits_class_meta_field_type_12_sub_class_id,
  input         io_class_meta_rsp_bits_class_meta_field_type_13_is_repeated,
  input  [4:0]  io_class_meta_rsp_bits_class_meta_field_type_13_field_type,
  input  [15:0] io_class_meta_rsp_bits_class_meta_field_type_13_sub_class_id,
  input         io_class_meta_rsp_bits_class_meta_field_type_14_is_repeated,
  input  [4:0]  io_class_meta_rsp_bits_class_meta_field_type_14_field_type,
  input  [15:0] io_class_meta_rsp_bits_class_meta_field_type_14_sub_class_id,
  input         io_class_meta_rsp_bits_class_meta_field_type_15_is_repeated,
  input  [4:0]  io_class_meta_rsp_bits_class_meta_field_type_15_field_type,
  input  [15:0] io_class_meta_rsp_bits_class_meta_field_type_15_sub_class_id,
  input         io_class_meta_rsp_bits_class_meta_field_type_16_is_repeated,
  input  [4:0]  io_class_meta_rsp_bits_class_meta_field_type_16_field_type,
  input  [15:0] io_class_meta_rsp_bits_class_meta_field_type_16_sub_class_id,
  input         io_class_meta_rsp_bits_class_meta_field_type_17_is_repeated,
  input  [4:0]  io_class_meta_rsp_bits_class_meta_field_type_17_field_type,
  input  [15:0] io_class_meta_rsp_bits_class_meta_field_type_17_sub_class_id,
  input         io_class_meta_rsp_bits_class_meta_field_type_18_is_repeated,
  input  [4:0]  io_class_meta_rsp_bits_class_meta_field_type_18_field_type,
  input  [15:0] io_class_meta_rsp_bits_class_meta_field_type_18_sub_class_id,
  input         io_class_meta_rsp_bits_class_meta_field_type_19_is_repeated,
  input  [4:0]  io_class_meta_rsp_bits_class_meta_field_type_19_field_type,
  input  [15:0] io_class_meta_rsp_bits_class_meta_field_type_19_sub_class_id,
  input         io_class_meta_rsp_bits_class_meta_field_type_20_is_repeated,
  input  [4:0]  io_class_meta_rsp_bits_class_meta_field_type_20_field_type,
  input  [15:0] io_class_meta_rsp_bits_class_meta_field_type_20_sub_class_id,
  input         io_class_meta_rsp_bits_class_meta_field_type_21_is_repeated,
  input  [4:0]  io_class_meta_rsp_bits_class_meta_field_type_21_field_type,
  input  [15:0] io_class_meta_rsp_bits_class_meta_field_type_21_sub_class_id,
  input         io_class_meta_rsp_bits_class_meta_field_type_22_is_repeated,
  input  [4:0]  io_class_meta_rsp_bits_class_meta_field_type_22_field_type,
  input  [15:0] io_class_meta_rsp_bits_class_meta_field_type_22_sub_class_id,
  input         io_class_meta_rsp_bits_class_meta_field_type_23_is_repeated,
  input  [4:0]  io_class_meta_rsp_bits_class_meta_field_type_23_field_type,
  input  [15:0] io_class_meta_rsp_bits_class_meta_field_type_23_sub_class_id,
  input         io_class_meta_rsp_bits_class_meta_field_type_24_is_repeated,
  input  [4:0]  io_class_meta_rsp_bits_class_meta_field_type_24_field_type,
  input  [15:0] io_class_meta_rsp_bits_class_meta_field_type_24_sub_class_id,
  input         io_class_meta_rsp_bits_class_meta_field_type_25_is_repeated,
  input  [4:0]  io_class_meta_rsp_bits_class_meta_field_type_25_field_type,
  input  [15:0] io_class_meta_rsp_bits_class_meta_field_type_25_sub_class_id,
  input         io_class_meta_rsp_bits_class_meta_field_type_26_is_repeated,
  input  [4:0]  io_class_meta_rsp_bits_class_meta_field_type_26_field_type,
  input  [15:0] io_class_meta_rsp_bits_class_meta_field_type_26_sub_class_id,
  input         io_class_meta_rsp_bits_class_meta_field_type_27_is_repeated,
  input  [4:0]  io_class_meta_rsp_bits_class_meta_field_type_27_field_type,
  input  [15:0] io_class_meta_rsp_bits_class_meta_field_type_27_sub_class_id,
  input         io_class_meta_rsp_bits_class_meta_field_type_28_is_repeated,
  input  [4:0]  io_class_meta_rsp_bits_class_meta_field_type_28_field_type,
  input  [15:0] io_class_meta_rsp_bits_class_meta_field_type_28_sub_class_id,
  input         io_class_meta_rsp_bits_class_meta_field_type_29_is_repeated,
  input  [4:0]  io_class_meta_rsp_bits_class_meta_field_type_29_field_type,
  input  [15:0] io_class_meta_rsp_bits_class_meta_field_type_29_sub_class_id,
  input         io_class_meta_rsp_bits_class_meta_field_type_30_is_repeated,
  input  [4:0]  io_class_meta_rsp_bits_class_meta_field_type_30_field_type,
  input  [15:0] io_class_meta_rsp_bits_class_meta_field_type_30_sub_class_id,
  input         io_class_meta_rsp_bits_class_meta_field_type_31_is_repeated,
  input  [4:0]  io_class_meta_rsp_bits_class_meta_field_type_31_field_type,
  input  [15:0] io_class_meta_rsp_bits_class_meta_field_type_31_sub_class_id,
  input         io_class_meta_rsp_bits_class_meta_field_type_32_is_repeated,
  input  [4:0]  io_class_meta_rsp_bits_class_meta_field_type_32_field_type,
  input  [15:0] io_class_meta_rsp_bits_class_meta_field_type_32_sub_class_id,
  input         io_done_ready,
  output        io_done_valid,
  output [31:0] counter_3_0,
  output [31:0] counter_2_0,
  output [31:0] counter_8,
  output [31:0] counter_1_1
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
  reg [31:0] _RAND_183;
  reg [31:0] _RAND_184;
  reg [31:0] _RAND_185;
  reg [31:0] _RAND_186;
  reg [31:0] _RAND_187;
  reg [31:0] _RAND_188;
  reg [31:0] _RAND_189;
  reg [31:0] _RAND_190;
  reg [31:0] _RAND_191;
  reg [31:0] _RAND_192;
  reg [31:0] _RAND_193;
  reg [31:0] _RAND_194;
  reg [31:0] _RAND_195;
  reg [31:0] _RAND_196;
  reg [31:0] _RAND_197;
  reg [31:0] _RAND_198;
  reg [31:0] _RAND_199;
  reg [31:0] _RAND_200;
  reg [31:0] _RAND_201;
  reg [31:0] _RAND_202;
  reg [31:0] _RAND_203;
  reg [31:0] _RAND_204;
  reg [31:0] _RAND_205;
  reg [31:0] _RAND_206;
  reg [31:0] _RAND_207;
  reg [31:0] _RAND_208;
  reg [31:0] _RAND_209;
  reg [31:0] _RAND_210;
  reg [31:0] _RAND_211;
  reg [31:0] _RAND_212;
  reg [31:0] _RAND_213;
  reg [31:0] _RAND_214;
  reg [31:0] _RAND_215;
  reg [31:0] _RAND_216;
  reg [31:0] _RAND_217;
  reg [31:0] _RAND_218;
  reg [31:0] _RAND_219;
  reg [31:0] _RAND_220;
  reg [31:0] _RAND_221;
  reg [31:0] _RAND_222;
  reg [31:0] _RAND_223;
  reg [31:0] _RAND_224;
  reg [31:0] _RAND_225;
  reg [31:0] _RAND_226;
  reg [31:0] _RAND_227;
  reg [31:0] _RAND_228;
  reg [31:0] _RAND_229;
  reg [31:0] _RAND_230;
  reg [31:0] _RAND_231;
  reg [31:0] _RAND_232;
  reg [31:0] _RAND_233;
  reg [31:0] _RAND_234;
  reg [31:0] _RAND_235;
  reg [31:0] _RAND_236;
  reg [31:0] _RAND_237;
  reg [31:0] _RAND_238;
  reg [31:0] _RAND_239;
  reg [31:0] _RAND_240;
  reg [31:0] _RAND_241;
  reg [31:0] _RAND_242;
  reg [31:0] _RAND_243;
  reg [31:0] _RAND_244;
  reg [31:0] _RAND_245;
  reg [31:0] _RAND_246;
  reg [31:0] _RAND_247;
  reg [31:0] _RAND_248;
  reg [31:0] _RAND_249;
  reg [31:0] _RAND_250;
  reg [31:0] _RAND_251;
  reg [31:0] _RAND_252;
  reg [31:0] _RAND_253;
  reg [31:0] _RAND_254;
  reg [31:0] _RAND_255;
  reg [31:0] _RAND_256;
  reg [31:0] _RAND_257;
  reg [31:0] _RAND_258;
  reg [31:0] _RAND_259;
  reg [31:0] _RAND_260;
  reg [31:0] _RAND_261;
  reg [31:0] _RAND_262;
  reg [31:0] _RAND_263;
  reg [31:0] _RAND_264;
  reg [31:0] _RAND_265;
  reg [31:0] _RAND_266;
  reg [31:0] _RAND_267;
  reg [31:0] _RAND_268;
  reg [31:0] _RAND_269;
  reg [31:0] _RAND_270;
  reg [31:0] _RAND_271;
  reg [31:0] _RAND_272;
  reg [31:0] _RAND_273;
  reg [31:0] _RAND_274;
  reg [31:0] _RAND_275;
  reg [31:0] _RAND_276;
  reg [31:0] _RAND_277;
  reg [31:0] _RAND_278;
  reg [31:0] _RAND_279;
  reg [31:0] _RAND_280;
  reg [31:0] _RAND_281;
  reg [31:0] _RAND_282;
  reg [31:0] _RAND_283;
  reg [31:0] _RAND_284;
  reg [31:0] _RAND_285;
  reg [31:0] _RAND_286;
  reg [31:0] _RAND_287;
  reg [31:0] _RAND_288;
  reg [31:0] _RAND_289;
  reg [31:0] _RAND_290;
  reg [31:0] _RAND_291;
  reg [31:0] _RAND_292;
  reg [31:0] _RAND_293;
  reg [31:0] _RAND_294;
  reg [31:0] _RAND_295;
  reg [31:0] _RAND_296;
  reg [31:0] _RAND_297;
  reg [31:0] _RAND_298;
  reg [31:0] _RAND_299;
  reg [31:0] _RAND_300;
  reg [31:0] _RAND_301;
  reg [31:0] _RAND_302;
  reg [31:0] _RAND_303;
  reg [31:0] _RAND_304;
  reg [31:0] _RAND_305;
  reg [31:0] _RAND_306;
  reg [31:0] _RAND_307;
  reg [31:0] _RAND_308;
  reg [31:0] _RAND_309;
  reg [31:0] _RAND_310;
  reg [31:0] _RAND_311;
  reg [31:0] _RAND_312;
  reg [31:0] _RAND_313;
  reg [31:0] _RAND_314;
  reg [31:0] _RAND_315;
  reg [31:0] _RAND_316;
  reg [31:0] _RAND_317;
  reg [31:0] _RAND_318;
  reg [31:0] _RAND_319;
  reg [31:0] _RAND_320;
  reg [31:0] _RAND_321;
  reg [31:0] _RAND_322;
  reg [31:0] _RAND_323;
  reg [31:0] _RAND_324;
  reg [31:0] _RAND_325;
  reg [31:0] _RAND_326;
  reg [31:0] _RAND_327;
  reg [31:0] _RAND_328;
  reg [31:0] _RAND_329;
  reg [31:0] _RAND_330;
  reg [31:0] _RAND_331;
  reg [31:0] _RAND_332;
  reg [31:0] _RAND_333;
  reg [31:0] _RAND_334;
  reg [31:0] _RAND_335;
  reg [31:0] _RAND_336;
  reg [31:0] _RAND_337;
  reg [31:0] _RAND_338;
  reg [31:0] _RAND_339;
  reg [31:0] _RAND_340;
  reg [31:0] _RAND_341;
  reg [31:0] _RAND_342;
  reg [31:0] _RAND_343;
  reg [31:0] _RAND_344;
  reg [31:0] _RAND_345;
  reg [31:0] _RAND_346;
  reg [31:0] _RAND_347;
  reg [31:0] _RAND_348;
  reg [31:0] _RAND_349;
  reg [31:0] _RAND_350;
  reg [31:0] _RAND_351;
  reg [31:0] _RAND_352;
  reg [31:0] _RAND_353;
  reg [31:0] _RAND_354;
  reg [31:0] _RAND_355;
  reg [31:0] _RAND_356;
  reg [31:0] _RAND_357;
  reg [31:0] _RAND_358;
  reg [31:0] _RAND_359;
  reg [31:0] _RAND_360;
  reg [31:0] _RAND_361;
  reg [31:0] _RAND_362;
  reg [31:0] _RAND_363;
  reg [31:0] _RAND_364;
  reg [31:0] _RAND_365;
  reg [31:0] _RAND_366;
  reg [31:0] _RAND_367;
  reg [31:0] _RAND_368;
  reg [31:0] _RAND_369;
  reg [31:0] _RAND_370;
  reg [31:0] _RAND_371;
  reg [31:0] _RAND_372;
  reg [31:0] _RAND_373;
  reg [31:0] _RAND_374;
  reg [31:0] _RAND_375;
  reg [31:0] _RAND_376;
  reg [31:0] _RAND_377;
  reg [31:0] _RAND_378;
  reg [31:0] _RAND_379;
  reg [31:0] _RAND_380;
  reg [31:0] _RAND_381;
  reg [31:0] _RAND_382;
  reg [31:0] _RAND_383;
  reg [31:0] _RAND_384;
  reg [31:0] _RAND_385;
  reg [31:0] _RAND_386;
  reg [31:0] _RAND_387;
  reg [31:0] _RAND_388;
  reg [31:0] _RAND_389;
  reg [31:0] _RAND_390;
  reg [31:0] _RAND_391;
  reg [31:0] _RAND_392;
  reg [31:0] _RAND_393;
  reg [31:0] _RAND_394;
  reg [31:0] _RAND_395;
  reg [31:0] _RAND_396;
  reg [31:0] _RAND_397;
  reg [31:0] _RAND_398;
  reg [31:0] _RAND_399;
  reg [31:0] _RAND_400;
  reg [31:0] _RAND_401;
  reg [31:0] _RAND_402;
  reg [31:0] _RAND_403;
  reg [31:0] _RAND_404;
  reg [31:0] _RAND_405;
  reg [31:0] _RAND_406;
  reg [31:0] _RAND_407;
  reg [31:0] _RAND_408;
  reg [31:0] _RAND_409;
  reg [31:0] _RAND_410;
  reg [31:0] _RAND_411;
  reg [31:0] _RAND_412;
  reg [31:0] _RAND_413;
  reg [31:0] _RAND_414;
  reg [31:0] _RAND_415;
  reg [31:0] _RAND_416;
  reg [31:0] _RAND_417;
  reg [31:0] _RAND_418;
  reg [31:0] _RAND_419;
  reg [31:0] _RAND_420;
  reg [31:0] _RAND_421;
  reg [31:0] _RAND_422;
  reg [31:0] _RAND_423;
  reg [31:0] _RAND_424;
  reg [31:0] _RAND_425;
  reg [31:0] _RAND_426;
  reg [31:0] _RAND_427;
  reg [31:0] _RAND_428;
  reg [31:0] _RAND_429;
  reg [31:0] _RAND_430;
  reg [31:0] _RAND_431;
  reg [31:0] _RAND_432;
  reg [31:0] _RAND_433;
  reg [31:0] _RAND_434;
  reg [31:0] _RAND_435;
  reg [31:0] _RAND_436;
  reg [31:0] _RAND_437;
  reg [31:0] _RAND_438;
  reg [31:0] _RAND_439;
  reg [31:0] _RAND_440;
  reg [31:0] _RAND_441;
  reg [31:0] _RAND_442;
  reg [31:0] _RAND_443;
  reg [31:0] _RAND_444;
  reg [31:0] _RAND_445;
  reg [31:0] _RAND_446;
  reg [31:0] _RAND_447;
  reg [31:0] _RAND_448;
  reg [31:0] _RAND_449;
  reg [31:0] _RAND_450;
  reg [31:0] _RAND_451;
  reg [31:0] _RAND_452;
  reg [31:0] _RAND_453;
  reg [31:0] _RAND_454;
  reg [31:0] _RAND_455;
  reg [31:0] _RAND_456;
  reg [31:0] _RAND_457;
  reg [31:0] _RAND_458;
  reg [31:0] _RAND_459;
  reg [31:0] _RAND_460;
  reg [31:0] _RAND_461;
  reg [31:0] _RAND_462;
  reg [31:0] _RAND_463;
  reg [31:0] _RAND_464;
  reg [31:0] _RAND_465;
  reg [31:0] _RAND_466;
  reg [31:0] _RAND_467;
  reg [31:0] _RAND_468;
  reg [31:0] _RAND_469;
  reg [31:0] _RAND_470;
  reg [31:0] _RAND_471;
  reg [31:0] _RAND_472;
  reg [31:0] _RAND_473;
  reg [31:0] _RAND_474;
  reg [31:0] _RAND_475;
  reg [31:0] _RAND_476;
  reg [31:0] _RAND_477;
  reg [31:0] _RAND_478;
  reg [31:0] _RAND_479;
  reg [31:0] _RAND_480;
  reg [31:0] _RAND_481;
  reg [31:0] _RAND_482;
  reg [31:0] _RAND_483;
  reg [31:0] _RAND_484;
  reg [31:0] _RAND_485;
  reg [31:0] _RAND_486;
  reg [31:0] _RAND_487;
  reg [31:0] _RAND_488;
  reg [31:0] _RAND_489;
  reg [31:0] _RAND_490;
  reg [31:0] _RAND_491;
  reg [31:0] _RAND_492;
  reg [31:0] _RAND_493;
  reg [31:0] _RAND_494;
  reg [31:0] _RAND_495;
  reg [31:0] _RAND_496;
  reg [31:0] _RAND_497;
  reg [31:0] _RAND_498;
  reg [31:0] _RAND_499;
  reg [31:0] _RAND_500;
  reg [31:0] _RAND_501;
  reg [31:0] _RAND_502;
  reg [31:0] _RAND_503;
  reg [31:0] _RAND_504;
  reg [31:0] _RAND_505;
  reg [31:0] _RAND_506;
  reg [31:0] _RAND_507;
  reg [31:0] _RAND_508;
  reg [31:0] _RAND_509;
  reg [31:0] _RAND_510;
  reg [31:0] _RAND_511;
  reg [31:0] _RAND_512;
  reg [31:0] _RAND_513;
  reg [31:0] _RAND_514;
  reg [31:0] _RAND_515;
  reg [31:0] _RAND_516;
  reg [31:0] _RAND_517;
  reg [31:0] _RAND_518;
  reg [31:0] _RAND_519;
  reg [31:0] _RAND_520;
  reg [31:0] _RAND_521;
  reg [31:0] _RAND_522;
  reg [31:0] _RAND_523;
  reg [31:0] _RAND_524;
  reg [31:0] _RAND_525;
  reg [31:0] _RAND_526;
  reg [31:0] _RAND_527;
  reg [31:0] _RAND_528;
  reg [31:0] _RAND_529;
  reg [31:0] _RAND_530;
  reg [31:0] _RAND_531;
  reg [31:0] _RAND_532;
  reg [31:0] _RAND_533;
  reg [31:0] _RAND_534;
  reg [31:0] _RAND_535;
  reg [31:0] _RAND_536;
  reg [31:0] _RAND_537;
  reg [31:0] _RAND_538;
  reg [31:0] _RAND_539;
  reg [31:0] _RAND_540;
  reg [31:0] _RAND_541;
  reg [31:0] _RAND_542;
  reg [31:0] _RAND_543;
  reg [31:0] _RAND_544;
  reg [31:0] _RAND_545;
  reg [31:0] _RAND_546;
  reg [31:0] _RAND_547;
  reg [31:0] _RAND_548;
  reg [31:0] _RAND_549;
  reg [31:0] _RAND_550;
  reg [31:0] _RAND_551;
  reg [31:0] _RAND_552;
  reg [31:0] _RAND_553;
  reg [31:0] _RAND_554;
  reg [31:0] _RAND_555;
  reg [31:0] _RAND_556;
  reg [31:0] _RAND_557;
  reg [31:0] _RAND_558;
  reg [31:0] _RAND_559;
  reg [31:0] _RAND_560;
  reg [31:0] _RAND_561;
  reg [31:0] _RAND_562;
  reg [31:0] _RAND_563;
  reg [31:0] _RAND_564;
  reg [31:0] _RAND_565;
  reg [31:0] _RAND_566;
  reg [31:0] _RAND_567;
  reg [31:0] _RAND_568;
  reg [31:0] _RAND_569;
  reg [31:0] _RAND_570;
  reg [31:0] _RAND_571;
  reg [31:0] _RAND_572;
  reg [31:0] _RAND_573;
  reg [31:0] _RAND_574;
  reg [31:0] _RAND_575;
  reg [31:0] _RAND_576;
  reg [31:0] _RAND_577;
  reg [31:0] _RAND_578;
  reg [31:0] _RAND_579;
  reg [31:0] _RAND_580;
  reg [31:0] _RAND_581;
  reg [31:0] _RAND_582;
  reg [31:0] _RAND_583;
  reg [31:0] _RAND_584;
  reg [31:0] _RAND_585;
  reg [31:0] _RAND_586;
  reg [31:0] _RAND_587;
  reg [31:0] _RAND_588;
  reg [31:0] _RAND_589;
  reg [31:0] _RAND_590;
  reg [31:0] _RAND_591;
  reg [31:0] _RAND_592;
  reg [31:0] _RAND_593;
  reg [31:0] _RAND_594;
  reg [31:0] _RAND_595;
  reg [31:0] _RAND_596;
  reg [31:0] _RAND_597;
  reg [31:0] _RAND_598;
  reg [31:0] _RAND_599;
  reg [31:0] _RAND_600;
  reg [31:0] _RAND_601;
  reg [31:0] _RAND_602;
  reg [31:0] _RAND_603;
  reg [31:0] _RAND_604;
  reg [31:0] _RAND_605;
  reg [31:0] _RAND_606;
  reg [31:0] _RAND_607;
  reg [31:0] _RAND_608;
  reg [31:0] _RAND_609;
  reg [31:0] _RAND_610;
  reg [31:0] _RAND_611;
  reg [31:0] _RAND_612;
  reg [31:0] _RAND_613;
  reg [31:0] _RAND_614;
  reg [31:0] _RAND_615;
  reg [31:0] _RAND_616;
  reg [31:0] _RAND_617;
  reg [31:0] _RAND_618;
  reg [31:0] _RAND_619;
  reg [31:0] _RAND_620;
  reg [31:0] _RAND_621;
  reg [31:0] _RAND_622;
  reg [31:0] _RAND_623;
  reg [31:0] _RAND_624;
  reg [31:0] _RAND_625;
  reg [31:0] _RAND_626;
  reg [31:0] _RAND_627;
  reg [31:0] _RAND_628;
  reg [31:0] _RAND_629;
  reg [31:0] _RAND_630;
  reg [31:0] _RAND_631;
  reg [31:0] _RAND_632;
  reg [31:0] _RAND_633;
  reg [31:0] _RAND_634;
  reg [31:0] _RAND_635;
  reg [31:0] _RAND_636;
  reg [31:0] _RAND_637;
  reg [31:0] _RAND_638;
  reg [31:0] _RAND_639;
  reg [31:0] _RAND_640;
  reg [31:0] _RAND_641;
  reg [31:0] _RAND_642;
  reg [31:0] _RAND_643;
  reg [31:0] _RAND_644;
  reg [31:0] _RAND_645;
  reg [31:0] _RAND_646;
  reg [31:0] _RAND_647;
  reg [31:0] _RAND_648;
  reg [31:0] _RAND_649;
  reg [31:0] _RAND_650;
  reg [31:0] _RAND_651;
  reg [31:0] _RAND_652;
  reg [31:0] _RAND_653;
  reg [31:0] _RAND_654;
  reg [31:0] _RAND_655;
  reg [31:0] _RAND_656;
  reg [31:0] _RAND_657;
  reg [31:0] _RAND_658;
  reg [31:0] _RAND_659;
  reg [31:0] _RAND_660;
  reg [31:0] _RAND_661;
  reg [31:0] _RAND_662;
  reg [31:0] _RAND_663;
  reg [31:0] _RAND_664;
  reg [31:0] _RAND_665;
  reg [31:0] _RAND_666;
  reg [31:0] _RAND_667;
  reg [31:0] _RAND_668;
  reg [31:0] _RAND_669;
  reg [31:0] _RAND_670;
  reg [31:0] _RAND_671;
  reg [31:0] _RAND_672;
  reg [31:0] _RAND_673;
  reg [31:0] _RAND_674;
  reg [31:0] _RAND_675;
  reg [31:0] _RAND_676;
  reg [31:0] _RAND_677;
  reg [31:0] _RAND_678;
  reg [31:0] _RAND_679;
  reg [31:0] _RAND_680;
  reg [31:0] _RAND_681;
  reg [31:0] _RAND_682;
  reg [31:0] _RAND_683;
  reg [31:0] _RAND_684;
  reg [31:0] _RAND_685;
  reg [31:0] _RAND_686;
  reg [31:0] _RAND_687;
  reg [31:0] _RAND_688;
  reg [31:0] _RAND_689;
  reg [31:0] _RAND_690;
  reg [31:0] _RAND_691;
  reg [31:0] _RAND_692;
  reg [31:0] _RAND_693;
  reg [31:0] _RAND_694;
  reg [31:0] _RAND_695;
  reg [31:0] _RAND_696;
  reg [31:0] _RAND_697;
  reg [31:0] _RAND_698;
  reg [31:0] _RAND_699;
  reg [31:0] _RAND_700;
  reg [31:0] _RAND_701;
  reg [31:0] _RAND_702;
  reg [31:0] _RAND_703;
  reg [31:0] _RAND_704;
  reg [31:0] _RAND_705;
  reg [31:0] _RAND_706;
  reg [31:0] _RAND_707;
  reg [31:0] _RAND_708;
  reg [31:0] _RAND_709;
  reg [31:0] _RAND_710;
  reg [31:0] _RAND_711;
  reg [31:0] _RAND_712;
  reg [31:0] _RAND_713;
  reg [31:0] _RAND_714;
  reg [31:0] _RAND_715;
  reg [31:0] _RAND_716;
  reg [31:0] _RAND_717;
  reg [31:0] _RAND_718;
  reg [31:0] _RAND_719;
  reg [31:0] _RAND_720;
  reg [31:0] _RAND_721;
  reg [31:0] _RAND_722;
  reg [31:0] _RAND_723;
  reg [31:0] _RAND_724;
  reg [31:0] _RAND_725;
  reg [31:0] _RAND_726;
  reg [31:0] _RAND_727;
  reg [31:0] _RAND_728;
  reg [31:0] _RAND_729;
  reg [31:0] _RAND_730;
  reg [31:0] _RAND_731;
  reg [31:0] _RAND_732;
  reg [31:0] _RAND_733;
  reg [31:0] _RAND_734;
  reg [31:0] _RAND_735;
  reg [31:0] _RAND_736;
  reg [31:0] _RAND_737;
  reg [31:0] _RAND_738;
  reg [31:0] _RAND_739;
  reg [31:0] _RAND_740;
  reg [31:0] _RAND_741;
  reg [31:0] _RAND_742;
  reg [31:0] _RAND_743;
  reg [31:0] _RAND_744;
  reg [31:0] _RAND_745;
  reg [31:0] _RAND_746;
  reg [31:0] _RAND_747;
  reg [31:0] _RAND_748;
  reg [31:0] _RAND_749;
  reg [31:0] _RAND_750;
  reg [31:0] _RAND_751;
  reg [31:0] _RAND_752;
  reg [31:0] _RAND_753;
  reg [31:0] _RAND_754;
  reg [31:0] _RAND_755;
  reg [31:0] _RAND_756;
  reg [31:0] _RAND_757;
  reg [31:0] _RAND_758;
  reg [31:0] _RAND_759;
  reg [31:0] _RAND_760;
  reg [31:0] _RAND_761;
  reg [31:0] _RAND_762;
  reg [31:0] _RAND_763;
  reg [31:0] _RAND_764;
  reg [31:0] _RAND_765;
  reg [31:0] _RAND_766;
  reg [31:0] _RAND_767;
  reg [31:0] _RAND_768;
  reg [31:0] _RAND_769;
  reg [31:0] _RAND_770;
  reg [31:0] _RAND_771;
  reg [31:0] _RAND_772;
  reg [31:0] _RAND_773;
  reg [31:0] _RAND_774;
  reg [31:0] _RAND_775;
  reg [31:0] _RAND_776;
  reg [31:0] _RAND_777;
  reg [31:0] _RAND_778;
  reg [31:0] _RAND_779;
  reg [31:0] _RAND_780;
  reg [31:0] _RAND_781;
  reg [31:0] _RAND_782;
  reg [31:0] _RAND_783;
  reg [31:0] _RAND_784;
  reg [31:0] _RAND_785;
  reg [31:0] _RAND_786;
  reg [31:0] _RAND_787;
  reg [31:0] _RAND_788;
  reg [31:0] _RAND_789;
  reg [31:0] _RAND_790;
  reg [31:0] _RAND_791;
  reg [31:0] _RAND_792;
  reg [31:0] _RAND_793;
  reg [31:0] _RAND_794;
  reg [31:0] _RAND_795;
  reg [31:0] _RAND_796;
  reg [31:0] _RAND_797;
  reg [31:0] _RAND_798;
  reg [31:0] _RAND_799;
  reg [31:0] _RAND_800;
  reg [31:0] _RAND_801;
  reg [31:0] _RAND_802;
  reg [31:0] _RAND_803;
  reg [31:0] _RAND_804;
  reg [31:0] _RAND_805;
  reg [31:0] _RAND_806;
  reg [31:0] _RAND_807;
  reg [31:0] _RAND_808;
  reg [31:0] _RAND_809;
  reg [31:0] _RAND_810;
  reg [31:0] _RAND_811;
  reg [31:0] _RAND_812;
  reg [31:0] _RAND_813;
  reg [31:0] _RAND_814;
  reg [31:0] _RAND_815;
  reg [31:0] _RAND_816;
  reg [31:0] _RAND_817;
  reg [31:0] _RAND_818;
  reg [31:0] _RAND_819;
  reg [31:0] _RAND_820;
  reg [31:0] _RAND_821;
  reg [31:0] _RAND_822;
  reg [31:0] _RAND_823;
  reg [31:0] _RAND_824;
  reg [31:0] _RAND_825;
  reg [31:0] _RAND_826;
  reg [31:0] _RAND_827;
  reg [31:0] _RAND_828;
  reg [31:0] _RAND_829;
  reg [31:0] _RAND_830;
  reg [31:0] _RAND_831;
  reg [31:0] _RAND_832;
  reg [31:0] _RAND_833;
  reg [31:0] _RAND_834;
  reg [31:0] _RAND_835;
  reg [31:0] _RAND_836;
  reg [31:0] _RAND_837;
  reg [31:0] _RAND_838;
  reg [31:0] _RAND_839;
  reg [31:0] _RAND_840;
  reg [31:0] _RAND_841;
  reg [31:0] _RAND_842;
  reg [31:0] _RAND_843;
  reg [31:0] _RAND_844;
  reg [31:0] _RAND_845;
  reg [31:0] _RAND_846;
  reg [31:0] _RAND_847;
  reg [31:0] _RAND_848;
  reg [31:0] _RAND_849;
  reg [31:0] _RAND_850;
  reg [31:0] _RAND_851;
  reg [31:0] _RAND_852;
  reg [31:0] _RAND_853;
  reg [31:0] _RAND_854;
  reg [31:0] _RAND_855;
  reg [31:0] _RAND_856;
  reg [31:0] _RAND_857;
  reg [31:0] _RAND_858;
  reg [31:0] _RAND_859;
  reg [31:0] _RAND_860;
  reg [31:0] _RAND_861;
  reg [31:0] _RAND_862;
  reg [31:0] _RAND_863;
  reg [31:0] _RAND_864;
  reg [31:0] _RAND_865;
  reg [31:0] _RAND_866;
  reg [31:0] _RAND_867;
  reg [31:0] _RAND_868;
  reg [31:0] _RAND_869;
  reg [31:0] _RAND_870;
  reg [31:0] _RAND_871;
  reg [31:0] _RAND_872;
  reg [31:0] _RAND_873;
  reg [31:0] _RAND_874;
  reg [31:0] _RAND_875;
  reg [31:0] _RAND_876;
  reg [31:0] _RAND_877;
  reg [31:0] _RAND_878;
  reg [31:0] _RAND_879;
  reg [31:0] _RAND_880;
  reg [31:0] _RAND_881;
  reg [31:0] _RAND_882;
  reg [31:0] _RAND_883;
  reg [31:0] _RAND_884;
  reg [31:0] _RAND_885;
  reg [31:0] _RAND_886;
  reg [31:0] _RAND_887;
  reg [31:0] _RAND_888;
  reg [31:0] _RAND_889;
  reg [31:0] _RAND_890;
  reg [31:0] _RAND_891;
  reg [31:0] _RAND_892;
  reg [31:0] _RAND_893;
  reg [31:0] _RAND_894;
  reg [31:0] _RAND_895;
  reg [31:0] _RAND_896;
  reg [31:0] _RAND_897;
  reg [31:0] _RAND_898;
  reg [31:0] _RAND_899;
  reg [31:0] _RAND_900;
  reg [31:0] _RAND_901;
  reg [31:0] _RAND_902;
  reg [31:0] _RAND_903;
  reg [31:0] _RAND_904;
  reg [31:0] _RAND_905;
  reg [31:0] _RAND_906;
  reg [31:0] _RAND_907;
  reg [31:0] _RAND_908;
  reg [31:0] _RAND_909;
  reg [31:0] _RAND_910;
  reg [31:0] _RAND_911;
  reg [31:0] _RAND_912;
  reg [31:0] _RAND_913;
  reg [31:0] _RAND_914;
  reg [31:0] _RAND_915;
  reg [31:0] _RAND_916;
  reg [31:0] _RAND_917;
  reg [31:0] _RAND_918;
  reg [31:0] _RAND_919;
  reg [31:0] _RAND_920;
  reg [31:0] _RAND_921;
  reg [31:0] _RAND_922;
  reg [31:0] _RAND_923;
  reg [31:0] _RAND_924;
  reg [31:0] _RAND_925;
  reg [31:0] _RAND_926;
  reg [31:0] _RAND_927;
  reg [31:0] _RAND_928;
  reg [31:0] _RAND_929;
  reg [31:0] _RAND_930;
  reg [31:0] _RAND_931;
  reg [31:0] _RAND_932;
  reg [31:0] _RAND_933;
  reg [31:0] _RAND_934;
  reg [31:0] _RAND_935;
  reg [31:0] _RAND_936;
  reg [31:0] _RAND_937;
  reg [31:0] _RAND_938;
  reg [31:0] _RAND_939;
  reg [31:0] _RAND_940;
  reg [31:0] _RAND_941;
  reg [31:0] _RAND_942;
  reg [31:0] _RAND_943;
  reg [31:0] _RAND_944;
  reg [31:0] _RAND_945;
  reg [31:0] _RAND_946;
  reg [31:0] _RAND_947;
  reg [31:0] _RAND_948;
  reg [31:0] _RAND_949;
  reg [31:0] _RAND_950;
  reg [31:0] _RAND_951;
  reg [31:0] _RAND_952;
  reg [31:0] _RAND_953;
  reg [31:0] _RAND_954;
  reg [31:0] _RAND_955;
  reg [31:0] _RAND_956;
  reg [31:0] _RAND_957;
  reg [31:0] _RAND_958;
  reg [31:0] _RAND_959;
  reg [31:0] _RAND_960;
  reg [31:0] _RAND_961;
  reg [31:0] _RAND_962;
  reg [31:0] _RAND_963;
  reg [31:0] _RAND_964;
  reg [31:0] _RAND_965;
  reg [31:0] _RAND_966;
  reg [31:0] _RAND_967;
  reg [31:0] _RAND_968;
  reg [31:0] _RAND_969;
  reg [31:0] _RAND_970;
  reg [31:0] _RAND_971;
  reg [31:0] _RAND_972;
  reg [31:0] _RAND_973;
  reg [31:0] _RAND_974;
  reg [31:0] _RAND_975;
  reg [31:0] _RAND_976;
  reg [31:0] _RAND_977;
  reg [31:0] _RAND_978;
  reg [31:0] _RAND_979;
  reg [31:0] _RAND_980;
  reg [31:0] _RAND_981;
  reg [31:0] _RAND_982;
  reg [31:0] _RAND_983;
  reg [31:0] _RAND_984;
  reg [31:0] _RAND_985;
  reg [31:0] _RAND_986;
  reg [31:0] _RAND_987;
  reg [31:0] _RAND_988;
  reg [31:0] _RAND_989;
  reg [31:0] _RAND_990;
  reg [31:0] _RAND_991;
  reg [31:0] _RAND_992;
  reg [31:0] _RAND_993;
  reg [31:0] _RAND_994;
  reg [31:0] _RAND_995;
  reg [31:0] _RAND_996;
  reg [31:0] _RAND_997;
  reg [31:0] _RAND_998;
  reg [31:0] _RAND_999;
  reg [31:0] _RAND_1000;
  reg [31:0] _RAND_1001;
  reg [31:0] _RAND_1002;
  reg [31:0] _RAND_1003;
  reg [31:0] _RAND_1004;
  reg [31:0] _RAND_1005;
  reg [31:0] _RAND_1006;
  reg [31:0] _RAND_1007;
  reg [31:0] _RAND_1008;
  reg [31:0] _RAND_1009;
  reg [31:0] _RAND_1010;
  reg [31:0] _RAND_1011;
  reg [31:0] _RAND_1012;
  reg [31:0] _RAND_1013;
  reg [31:0] _RAND_1014;
  reg [31:0] _RAND_1015;
  reg [31:0] _RAND_1016;
  reg [31:0] _RAND_1017;
  reg [31:0] _RAND_1018;
  reg [31:0] _RAND_1019;
  reg [31:0] _RAND_1020;
  reg [31:0] _RAND_1021;
  reg [31:0] _RAND_1022;
  reg [31:0] _RAND_1023;
  reg [31:0] _RAND_1024;
  reg [31:0] _RAND_1025;
  reg [31:0] _RAND_1026;
  reg [31:0] _RAND_1027;
  reg [31:0] _RAND_1028;
  reg [31:0] _RAND_1029;
  reg [31:0] _RAND_1030;
  reg [31:0] _RAND_1031;
  reg [31:0] _RAND_1032;
  reg [31:0] _RAND_1033;
  reg [31:0] _RAND_1034;
  reg [31:0] _RAND_1035;
  reg [31:0] _RAND_1036;
  reg [31:0] _RAND_1037;
  reg [31:0] _RAND_1038;
  reg [31:0] _RAND_1039;
  reg [31:0] _RAND_1040;
  reg [31:0] _RAND_1041;
  reg [31:0] _RAND_1042;
  reg [31:0] _RAND_1043;
  reg [31:0] _RAND_1044;
  reg [31:0] _RAND_1045;
  reg [31:0] _RAND_1046;
  reg [31:0] _RAND_1047;
  reg [31:0] _RAND_1048;
  reg [31:0] _RAND_1049;
  reg [31:0] _RAND_1050;
  reg [31:0] _RAND_1051;
  reg [31:0] _RAND_1052;
  reg [31:0] _RAND_1053;
  reg [31:0] _RAND_1054;
  reg [31:0] _RAND_1055;
  reg [31:0] _RAND_1056;
  reg [31:0] _RAND_1057;
  reg [31:0] _RAND_1058;
  reg [31:0] _RAND_1059;
  reg [31:0] _RAND_1060;
  reg [31:0] _RAND_1061;
  reg [31:0] _RAND_1062;
  reg [31:0] _RAND_1063;
  reg [31:0] _RAND_1064;
  reg [31:0] _RAND_1065;
  reg [31:0] _RAND_1066;
  reg [31:0] _RAND_1067;
  reg [31:0] _RAND_1068;
  reg [31:0] _RAND_1069;
  reg [31:0] _RAND_1070;
  reg [31:0] _RAND_1071;
  reg [31:0] _RAND_1072;
  reg [31:0] _RAND_1073;
  reg [31:0] _RAND_1074;
  reg [31:0] _RAND_1075;
  reg [31:0] _RAND_1076;
  reg [31:0] _RAND_1077;
  reg [31:0] _RAND_1078;
  reg [31:0] _RAND_1079;
  reg [31:0] _RAND_1080;
  reg [31:0] _RAND_1081;
  reg [31:0] _RAND_1082;
  reg [31:0] _RAND_1083;
  reg [31:0] _RAND_1084;
  reg [31:0] _RAND_1085;
  reg [31:0] _RAND_1086;
  reg [31:0] _RAND_1087;
  reg [31:0] _RAND_1088;
  reg [31:0] _RAND_1089;
  reg [31:0] _RAND_1090;
  reg [31:0] _RAND_1091;
  reg [31:0] _RAND_1092;
  reg [31:0] _RAND_1093;
  reg [31:0] _RAND_1094;
  reg [31:0] _RAND_1095;
  reg [31:0] _RAND_1096;
  reg [31:0] _RAND_1097;
  reg [31:0] _RAND_1098;
  reg [31:0] _RAND_1099;
  reg [31:0] _RAND_1100;
  reg [31:0] _RAND_1101;
  reg [31:0] _RAND_1102;
  reg [31:0] _RAND_1103;
  reg [31:0] _RAND_1104;
  reg [31:0] _RAND_1105;
  reg [31:0] _RAND_1106;
  reg [31:0] _RAND_1107;
  reg [31:0] _RAND_1108;
  reg [31:0] _RAND_1109;
  reg [31:0] _RAND_1110;
  reg [31:0] _RAND_1111;
  reg [31:0] _RAND_1112;
  reg [31:0] _RAND_1113;
  reg [31:0] _RAND_1114;
  reg [31:0] _RAND_1115;
  reg [31:0] _RAND_1116;
  reg [31:0] _RAND_1117;
  reg [31:0] _RAND_1118;
  reg [31:0] _RAND_1119;
  reg [31:0] _RAND_1120;
  reg [31:0] _RAND_1121;
  reg [31:0] _RAND_1122;
  reg [31:0] _RAND_1123;
  reg [31:0] _RAND_1124;
  reg [31:0] _RAND_1125;
  reg [31:0] _RAND_1126;
  reg [31:0] _RAND_1127;
  reg [31:0] _RAND_1128;
  reg [31:0] _RAND_1129;
  reg [31:0] _RAND_1130;
  reg [31:0] _RAND_1131;
  reg [31:0] _RAND_1132;
  reg [31:0] _RAND_1133;
  reg [31:0] _RAND_1134;
  reg [31:0] _RAND_1135;
  reg [31:0] _RAND_1136;
  reg [31:0] _RAND_1137;
  reg [31:0] _RAND_1138;
  reg [31:0] _RAND_1139;
  reg [31:0] _RAND_1140;
  reg [31:0] _RAND_1141;
  reg [31:0] _RAND_1142;
  reg [31:0] _RAND_1143;
  reg [31:0] _RAND_1144;
  reg [31:0] _RAND_1145;
  reg [31:0] _RAND_1146;
  reg [31:0] _RAND_1147;
  reg [31:0] _RAND_1148;
  reg [31:0] _RAND_1149;
  reg [31:0] _RAND_1150;
  reg [31:0] _RAND_1151;
  reg [31:0] _RAND_1152;
  reg [31:0] _RAND_1153;
  reg [31:0] _RAND_1154;
  reg [31:0] _RAND_1155;
  reg [31:0] _RAND_1156;
  reg [31:0] _RAND_1157;
  reg [31:0] _RAND_1158;
  reg [31:0] _RAND_1159;
  reg [31:0] _RAND_1160;
  reg [31:0] _RAND_1161;
  reg [31:0] _RAND_1162;
  reg [31:0] _RAND_1163;
  reg [31:0] _RAND_1164;
  reg [31:0] _RAND_1165;
  reg [31:0] _RAND_1166;
  reg [31:0] _RAND_1167;
  reg [31:0] _RAND_1168;
  reg [31:0] _RAND_1169;
  reg [31:0] _RAND_1170;
  reg [31:0] _RAND_1171;
  reg [31:0] _RAND_1172;
  reg [31:0] _RAND_1173;
  reg [31:0] _RAND_1174;
  reg [31:0] _RAND_1175;
  reg [31:0] _RAND_1176;
  reg [31:0] _RAND_1177;
  reg [31:0] _RAND_1178;
  reg [31:0] _RAND_1179;
  reg [31:0] _RAND_1180;
  reg [31:0] _RAND_1181;
  reg [31:0] _RAND_1182;
  reg [31:0] _RAND_1183;
  reg [31:0] _RAND_1184;
  reg [31:0] _RAND_1185;
  reg [31:0] _RAND_1186;
  reg [31:0] _RAND_1187;
  reg [31:0] _RAND_1188;
  reg [31:0] _RAND_1189;
  reg [31:0] _RAND_1190;
  reg [31:0] _RAND_1191;
  reg [31:0] _RAND_1192;
  reg [31:0] _RAND_1193;
  reg [31:0] _RAND_1194;
  reg [31:0] _RAND_1195;
  reg [31:0] _RAND_1196;
  reg [31:0] _RAND_1197;
  reg [31:0] _RAND_1198;
  reg [31:0] _RAND_1199;
  reg [31:0] _RAND_1200;
  reg [31:0] _RAND_1201;
  reg [31:0] _RAND_1202;
  reg [31:0] _RAND_1203;
  reg [31:0] _RAND_1204;
  reg [31:0] _RAND_1205;
  reg [31:0] _RAND_1206;
  reg [31:0] _RAND_1207;
  reg [31:0] _RAND_1208;
  reg [31:0] _RAND_1209;
  reg [31:0] _RAND_1210;
  reg [31:0] _RAND_1211;
  reg [31:0] _RAND_1212;
  reg [31:0] _RAND_1213;
  reg [31:0] _RAND_1214;
  reg [31:0] _RAND_1215;
  reg [31:0] _RAND_1216;
  reg [31:0] _RAND_1217;
  reg [31:0] _RAND_1218;
  reg [31:0] _RAND_1219;
  reg [31:0] _RAND_1220;
  reg [31:0] _RAND_1221;
  reg [31:0] _RAND_1222;
  reg [31:0] _RAND_1223;
  reg [31:0] _RAND_1224;
  reg [31:0] _RAND_1225;
  reg [31:0] _RAND_1226;
  reg [31:0] _RAND_1227;
  reg [31:0] _RAND_1228;
  reg [31:0] _RAND_1229;
  reg [31:0] _RAND_1230;
  reg [31:0] _RAND_1231;
  reg [31:0] _RAND_1232;
  reg [31:0] _RAND_1233;
  reg [31:0] _RAND_1234;
  reg [31:0] _RAND_1235;
  reg [31:0] _RAND_1236;
  reg [31:0] _RAND_1237;
  reg [31:0] _RAND_1238;
  reg [31:0] _RAND_1239;
  reg [31:0] _RAND_1240;
  reg [31:0] _RAND_1241;
  reg [31:0] _RAND_1242;
  reg [31:0] _RAND_1243;
  reg [31:0] _RAND_1244;
  reg [31:0] _RAND_1245;
  reg [31:0] _RAND_1246;
  reg [31:0] _RAND_1247;
  reg [31:0] _RAND_1248;
  reg [31:0] _RAND_1249;
  reg [31:0] _RAND_1250;
  reg [31:0] _RAND_1251;
  reg [31:0] _RAND_1252;
  reg [31:0] _RAND_1253;
  reg [31:0] _RAND_1254;
  reg [31:0] _RAND_1255;
  reg [31:0] _RAND_1256;
  reg [31:0] _RAND_1257;
  reg [31:0] _RAND_1258;
  reg [31:0] _RAND_1259;
  reg [31:0] _RAND_1260;
  reg [31:0] _RAND_1261;
  reg [31:0] _RAND_1262;
  reg [31:0] _RAND_1263;
  reg [31:0] _RAND_1264;
  reg [31:0] _RAND_1265;
  reg [31:0] _RAND_1266;
  reg [31:0] _RAND_1267;
  reg [31:0] _RAND_1268;
  reg [31:0] _RAND_1269;
  reg [31:0] _RAND_1270;
  reg [31:0] _RAND_1271;
  reg [31:0] _RAND_1272;
  reg [31:0] _RAND_1273;
  reg [31:0] _RAND_1274;
  reg [31:0] _RAND_1275;
  reg [31:0] _RAND_1276;
  reg [31:0] _RAND_1277;
  reg [31:0] _RAND_1278;
  reg [31:0] _RAND_1279;
  reg [31:0] _RAND_1280;
  reg [31:0] _RAND_1281;
  reg [31:0] _RAND_1282;
  reg [31:0] _RAND_1283;
  reg [31:0] _RAND_1284;
  reg [31:0] _RAND_1285;
  reg [31:0] _RAND_1286;
  reg [31:0] _RAND_1287;
  reg [31:0] _RAND_1288;
  reg [31:0] _RAND_1289;
  reg [31:0] _RAND_1290;
  reg [31:0] _RAND_1291;
  reg [31:0] _RAND_1292;
  reg [31:0] _RAND_1293;
  reg [31:0] _RAND_1294;
  reg [31:0] _RAND_1295;
  reg [31:0] _RAND_1296;
  reg [31:0] _RAND_1297;
  reg [31:0] _RAND_1298;
  reg [31:0] _RAND_1299;
  reg [31:0] _RAND_1300;
  reg [31:0] _RAND_1301;
  reg [31:0] _RAND_1302;
  reg [31:0] _RAND_1303;
  reg [31:0] _RAND_1304;
  reg [31:0] _RAND_1305;
  reg [31:0] _RAND_1306;
  reg [31:0] _RAND_1307;
  reg [31:0] _RAND_1308;
  reg [31:0] _RAND_1309;
  reg [31:0] _RAND_1310;
  reg [31:0] _RAND_1311;
  reg [31:0] _RAND_1312;
  reg [31:0] _RAND_1313;
  reg [31:0] _RAND_1314;
  reg [31:0] _RAND_1315;
  reg [31:0] _RAND_1316;
  reg [31:0] _RAND_1317;
  reg [31:0] _RAND_1318;
  reg [31:0] _RAND_1319;
  reg [31:0] _RAND_1320;
  reg [31:0] _RAND_1321;
  reg [31:0] _RAND_1322;
  reg [31:0] _RAND_1323;
  reg [31:0] _RAND_1324;
  reg [31:0] _RAND_1325;
  reg [31:0] _RAND_1326;
  reg [31:0] _RAND_1327;
  reg [31:0] _RAND_1328;
  reg [31:0] _RAND_1329;
  reg [31:0] _RAND_1330;
  reg [31:0] _RAND_1331;
  reg [31:0] _RAND_1332;
  reg [31:0] _RAND_1333;
  reg [31:0] _RAND_1334;
  reg [31:0] _RAND_1335;
  reg [31:0] _RAND_1336;
  reg [31:0] _RAND_1337;
  reg [31:0] _RAND_1338;
  reg [31:0] _RAND_1339;
  reg [31:0] _RAND_1340;
  reg [31:0] _RAND_1341;
  reg [31:0] _RAND_1342;
  reg [31:0] _RAND_1343;
  reg [31:0] _RAND_1344;
  reg [31:0] _RAND_1345;
  reg [31:0] _RAND_1346;
  reg [31:0] _RAND_1347;
  reg [31:0] _RAND_1348;
  reg [31:0] _RAND_1349;
  reg [31:0] _RAND_1350;
  reg [31:0] _RAND_1351;
  reg [31:0] _RAND_1352;
  reg [31:0] _RAND_1353;
  reg [31:0] _RAND_1354;
  reg [31:0] _RAND_1355;
  reg [31:0] _RAND_1356;
  reg [31:0] _RAND_1357;
  reg [31:0] _RAND_1358;
  reg [31:0] _RAND_1359;
  reg [31:0] _RAND_1360;
  reg [31:0] _RAND_1361;
  reg [31:0] _RAND_1362;
  reg [31:0] _RAND_1363;
  reg [31:0] _RAND_1364;
  reg [31:0] _RAND_1365;
  reg [31:0] _RAND_1366;
  reg [31:0] _RAND_1367;
  reg [31:0] _RAND_1368;
  reg [31:0] _RAND_1369;
  reg [31:0] _RAND_1370;
  reg [31:0] _RAND_1371;
  reg [31:0] _RAND_1372;
  reg [31:0] _RAND_1373;
  reg [31:0] _RAND_1374;
  reg [31:0] _RAND_1375;
  reg [31:0] _RAND_1376;
  reg [31:0] _RAND_1377;
  reg [31:0] _RAND_1378;
  reg [31:0] _RAND_1379;
  reg [31:0] _RAND_1380;
  reg [31:0] _RAND_1381;
  reg [31:0] _RAND_1382;
  reg [31:0] _RAND_1383;
  reg [31:0] _RAND_1384;
  reg [31:0] _RAND_1385;
  reg [31:0] _RAND_1386;
  reg [31:0] _RAND_1387;
  reg [31:0] _RAND_1388;
  reg [31:0] _RAND_1389;
  reg [31:0] _RAND_1390;
  reg [31:0] _RAND_1391;
  reg [31:0] _RAND_1392;
  reg [31:0] _RAND_1393;
  reg [31:0] _RAND_1394;
  reg [31:0] _RAND_1395;
  reg [31:0] _RAND_1396;
  reg [31:0] _RAND_1397;
  reg [31:0] _RAND_1398;
  reg [31:0] _RAND_1399;
  reg [31:0] _RAND_1400;
  reg [31:0] _RAND_1401;
  reg [31:0] _RAND_1402;
  reg [31:0] _RAND_1403;
  reg [31:0] _RAND_1404;
  reg [31:0] _RAND_1405;
  reg [31:0] _RAND_1406;
  reg [31:0] _RAND_1407;
  reg [31:0] _RAND_1408;
  reg [31:0] _RAND_1409;
  reg [31:0] _RAND_1410;
  reg [31:0] _RAND_1411;
  reg [31:0] _RAND_1412;
  reg [31:0] _RAND_1413;
  reg [31:0] _RAND_1414;
  reg [31:0] _RAND_1415;
  reg [31:0] _RAND_1416;
  reg [31:0] _RAND_1417;
  reg [31:0] _RAND_1418;
  reg [31:0] _RAND_1419;
  reg [31:0] _RAND_1420;
  reg [31:0] _RAND_1421;
  reg [31:0] _RAND_1422;
  reg [31:0] _RAND_1423;
  reg [31:0] _RAND_1424;
  reg [31:0] _RAND_1425;
  reg [31:0] _RAND_1426;
  reg [31:0] _RAND_1427;
  reg [31:0] _RAND_1428;
  reg [31:0] _RAND_1429;
  reg [31:0] _RAND_1430;
  reg [31:0] _RAND_1431;
  reg [31:0] _RAND_1432;
  reg [31:0] _RAND_1433;
  reg [31:0] _RAND_1434;
  reg [31:0] _RAND_1435;
  reg [31:0] _RAND_1436;
  reg [31:0] _RAND_1437;
  reg [31:0] _RAND_1438;
  reg [31:0] _RAND_1439;
  reg [31:0] _RAND_1440;
  reg [31:0] _RAND_1441;
  reg [31:0] _RAND_1442;
  reg [31:0] _RAND_1443;
  reg [31:0] _RAND_1444;
  reg [31:0] _RAND_1445;
  reg [31:0] _RAND_1446;
  reg [31:0] _RAND_1447;
  reg [31:0] _RAND_1448;
  reg [31:0] _RAND_1449;
  reg [31:0] _RAND_1450;
  reg [31:0] _RAND_1451;
  reg [31:0] _RAND_1452;
  reg [31:0] _RAND_1453;
  reg [31:0] _RAND_1454;
  reg [31:0] _RAND_1455;
  reg [31:0] _RAND_1456;
  reg [31:0] _RAND_1457;
  reg [31:0] _RAND_1458;
  reg [31:0] _RAND_1459;
  reg [31:0] _RAND_1460;
  reg [31:0] _RAND_1461;
  reg [31:0] _RAND_1462;
  reg [31:0] _RAND_1463;
  reg [31:0] _RAND_1464;
  reg [31:0] _RAND_1465;
  reg [31:0] _RAND_1466;
  reg [31:0] _RAND_1467;
  reg [31:0] _RAND_1468;
  reg [31:0] _RAND_1469;
  reg [31:0] _RAND_1470;
  reg [31:0] _RAND_1471;
  reg [31:0] _RAND_1472;
  reg [31:0] _RAND_1473;
  reg [31:0] _RAND_1474;
  reg [31:0] _RAND_1475;
  reg [31:0] _RAND_1476;
  reg [31:0] _RAND_1477;
  reg [31:0] _RAND_1478;
  reg [31:0] _RAND_1479;
  reg [31:0] _RAND_1480;
  reg [31:0] _RAND_1481;
  reg [31:0] _RAND_1482;
  reg [31:0] _RAND_1483;
  reg [31:0] _RAND_1484;
  reg [31:0] _RAND_1485;
  reg [31:0] _RAND_1486;
  reg [31:0] _RAND_1487;
  reg [31:0] _RAND_1488;
  reg [31:0] _RAND_1489;
  reg [31:0] _RAND_1490;
  reg [31:0] _RAND_1491;
  reg [31:0] _RAND_1492;
  reg [31:0] _RAND_1493;
  reg [31:0] _RAND_1494;
  reg [31:0] _RAND_1495;
  reg [31:0] _RAND_1496;
  reg [31:0] _RAND_1497;
  reg [31:0] _RAND_1498;
  reg [31:0] _RAND_1499;
  reg [31:0] _RAND_1500;
  reg [31:0] _RAND_1501;
  reg [31:0] _RAND_1502;
  reg [31:0] _RAND_1503;
  reg [31:0] _RAND_1504;
  reg [63:0] _RAND_1505;
  reg [31:0] _RAND_1506;
  reg [31:0] _RAND_1507;
  reg [31:0] _RAND_1508;
  reg [31:0] _RAND_1509;
  reg [31:0] _RAND_1510;
  reg [31:0] _RAND_1511;
  reg [31:0] _RAND_1512;
  reg [31:0] _RAND_1513;
`endif // RANDOMIZE_REG_INIT
  wire  meta_in_fifo_clock; // @[XQueue.scala 35:23]
  wire  meta_in_fifo_reset; // @[XQueue.scala 35:23]
  wire  meta_in_fifo_io_in_ready; // @[XQueue.scala 35:23]
  wire  meta_in_fifo_io_in_valid; // @[XQueue.scala 35:23]
  wire [9:0] meta_in_fifo_io_in_bits_class_id; // @[XQueue.scala 35:23]
  wire [63:0] meta_in_fifo_io_in_bits_host_base_addr; // @[XQueue.scala 35:23]
  wire  meta_in_fifo_io_out_ready; // @[XQueue.scala 35:23]
  wire  meta_in_fifo_io_out_valid; // @[XQueue.scala 35:23]
  wire [9:0] meta_in_fifo_io_out_bits_class_id; // @[XQueue.scala 35:23]
  wire [63:0] meta_in_fifo_io_out_bits_host_base_addr; // @[XQueue.scala 35:23]
  wire  class_meta_rsp_fifo_clock; // @[XQueue.scala 35:23]
  wire  class_meta_rsp_fifo_reset; // @[XQueue.scala 35:23]
  wire  class_meta_rsp_fifo_io_in_valid; // @[XQueue.scala 35:23]
  wire [7:0] class_meta_rsp_fifo_io_in_bits_class_meta_max_field_num; // @[XQueue.scala 35:23]
  wire  class_meta_rsp_fifo_io_in_bits_class_meta_field_type_0_is_repeated; // @[XQueue.scala 35:23]
  wire [4:0] class_meta_rsp_fifo_io_in_bits_class_meta_field_type_0_field_type; // @[XQueue.scala 35:23]
  wire [15:0] class_meta_rsp_fifo_io_in_bits_class_meta_field_type_0_sub_class_id; // @[XQueue.scala 35:23]
  wire  class_meta_rsp_fifo_io_in_bits_class_meta_field_type_1_is_repeated; // @[XQueue.scala 35:23]
  wire [4:0] class_meta_rsp_fifo_io_in_bits_class_meta_field_type_1_field_type; // @[XQueue.scala 35:23]
  wire [15:0] class_meta_rsp_fifo_io_in_bits_class_meta_field_type_1_sub_class_id; // @[XQueue.scala 35:23]
  wire  class_meta_rsp_fifo_io_in_bits_class_meta_field_type_2_is_repeated; // @[XQueue.scala 35:23]
  wire [4:0] class_meta_rsp_fifo_io_in_bits_class_meta_field_type_2_field_type; // @[XQueue.scala 35:23]
  wire [15:0] class_meta_rsp_fifo_io_in_bits_class_meta_field_type_2_sub_class_id; // @[XQueue.scala 35:23]
  wire  class_meta_rsp_fifo_io_in_bits_class_meta_field_type_3_is_repeated; // @[XQueue.scala 35:23]
  wire [4:0] class_meta_rsp_fifo_io_in_bits_class_meta_field_type_3_field_type; // @[XQueue.scala 35:23]
  wire [15:0] class_meta_rsp_fifo_io_in_bits_class_meta_field_type_3_sub_class_id; // @[XQueue.scala 35:23]
  wire  class_meta_rsp_fifo_io_in_bits_class_meta_field_type_4_is_repeated; // @[XQueue.scala 35:23]
  wire [4:0] class_meta_rsp_fifo_io_in_bits_class_meta_field_type_4_field_type; // @[XQueue.scala 35:23]
  wire [15:0] class_meta_rsp_fifo_io_in_bits_class_meta_field_type_4_sub_class_id; // @[XQueue.scala 35:23]
  wire  class_meta_rsp_fifo_io_in_bits_class_meta_field_type_5_is_repeated; // @[XQueue.scala 35:23]
  wire [4:0] class_meta_rsp_fifo_io_in_bits_class_meta_field_type_5_field_type; // @[XQueue.scala 35:23]
  wire [15:0] class_meta_rsp_fifo_io_in_bits_class_meta_field_type_5_sub_class_id; // @[XQueue.scala 35:23]
  wire  class_meta_rsp_fifo_io_in_bits_class_meta_field_type_6_is_repeated; // @[XQueue.scala 35:23]
  wire [4:0] class_meta_rsp_fifo_io_in_bits_class_meta_field_type_6_field_type; // @[XQueue.scala 35:23]
  wire [15:0] class_meta_rsp_fifo_io_in_bits_class_meta_field_type_6_sub_class_id; // @[XQueue.scala 35:23]
  wire  class_meta_rsp_fifo_io_in_bits_class_meta_field_type_7_is_repeated; // @[XQueue.scala 35:23]
  wire [4:0] class_meta_rsp_fifo_io_in_bits_class_meta_field_type_7_field_type; // @[XQueue.scala 35:23]
  wire [15:0] class_meta_rsp_fifo_io_in_bits_class_meta_field_type_7_sub_class_id; // @[XQueue.scala 35:23]
  wire  class_meta_rsp_fifo_io_in_bits_class_meta_field_type_8_is_repeated; // @[XQueue.scala 35:23]
  wire [4:0] class_meta_rsp_fifo_io_in_bits_class_meta_field_type_8_field_type; // @[XQueue.scala 35:23]
  wire [15:0] class_meta_rsp_fifo_io_in_bits_class_meta_field_type_8_sub_class_id; // @[XQueue.scala 35:23]
  wire  class_meta_rsp_fifo_io_in_bits_class_meta_field_type_9_is_repeated; // @[XQueue.scala 35:23]
  wire [4:0] class_meta_rsp_fifo_io_in_bits_class_meta_field_type_9_field_type; // @[XQueue.scala 35:23]
  wire [15:0] class_meta_rsp_fifo_io_in_bits_class_meta_field_type_9_sub_class_id; // @[XQueue.scala 35:23]
  wire  class_meta_rsp_fifo_io_in_bits_class_meta_field_type_10_is_repeated; // @[XQueue.scala 35:23]
  wire [4:0] class_meta_rsp_fifo_io_in_bits_class_meta_field_type_10_field_type; // @[XQueue.scala 35:23]
  wire [15:0] class_meta_rsp_fifo_io_in_bits_class_meta_field_type_10_sub_class_id; // @[XQueue.scala 35:23]
  wire  class_meta_rsp_fifo_io_in_bits_class_meta_field_type_11_is_repeated; // @[XQueue.scala 35:23]
  wire [4:0] class_meta_rsp_fifo_io_in_bits_class_meta_field_type_11_field_type; // @[XQueue.scala 35:23]
  wire [15:0] class_meta_rsp_fifo_io_in_bits_class_meta_field_type_11_sub_class_id; // @[XQueue.scala 35:23]
  wire  class_meta_rsp_fifo_io_in_bits_class_meta_field_type_12_is_repeated; // @[XQueue.scala 35:23]
  wire [4:0] class_meta_rsp_fifo_io_in_bits_class_meta_field_type_12_field_type; // @[XQueue.scala 35:23]
  wire [15:0] class_meta_rsp_fifo_io_in_bits_class_meta_field_type_12_sub_class_id; // @[XQueue.scala 35:23]
  wire  class_meta_rsp_fifo_io_in_bits_class_meta_field_type_13_is_repeated; // @[XQueue.scala 35:23]
  wire [4:0] class_meta_rsp_fifo_io_in_bits_class_meta_field_type_13_field_type; // @[XQueue.scala 35:23]
  wire [15:0] class_meta_rsp_fifo_io_in_bits_class_meta_field_type_13_sub_class_id; // @[XQueue.scala 35:23]
  wire  class_meta_rsp_fifo_io_in_bits_class_meta_field_type_14_is_repeated; // @[XQueue.scala 35:23]
  wire [4:0] class_meta_rsp_fifo_io_in_bits_class_meta_field_type_14_field_type; // @[XQueue.scala 35:23]
  wire [15:0] class_meta_rsp_fifo_io_in_bits_class_meta_field_type_14_sub_class_id; // @[XQueue.scala 35:23]
  wire  class_meta_rsp_fifo_io_in_bits_class_meta_field_type_15_is_repeated; // @[XQueue.scala 35:23]
  wire [4:0] class_meta_rsp_fifo_io_in_bits_class_meta_field_type_15_field_type; // @[XQueue.scala 35:23]
  wire [15:0] class_meta_rsp_fifo_io_in_bits_class_meta_field_type_15_sub_class_id; // @[XQueue.scala 35:23]
  wire  class_meta_rsp_fifo_io_in_bits_class_meta_field_type_16_is_repeated; // @[XQueue.scala 35:23]
  wire [4:0] class_meta_rsp_fifo_io_in_bits_class_meta_field_type_16_field_type; // @[XQueue.scala 35:23]
  wire [15:0] class_meta_rsp_fifo_io_in_bits_class_meta_field_type_16_sub_class_id; // @[XQueue.scala 35:23]
  wire  class_meta_rsp_fifo_io_in_bits_class_meta_field_type_17_is_repeated; // @[XQueue.scala 35:23]
  wire [4:0] class_meta_rsp_fifo_io_in_bits_class_meta_field_type_17_field_type; // @[XQueue.scala 35:23]
  wire [15:0] class_meta_rsp_fifo_io_in_bits_class_meta_field_type_17_sub_class_id; // @[XQueue.scala 35:23]
  wire  class_meta_rsp_fifo_io_in_bits_class_meta_field_type_18_is_repeated; // @[XQueue.scala 35:23]
  wire [4:0] class_meta_rsp_fifo_io_in_bits_class_meta_field_type_18_field_type; // @[XQueue.scala 35:23]
  wire [15:0] class_meta_rsp_fifo_io_in_bits_class_meta_field_type_18_sub_class_id; // @[XQueue.scala 35:23]
  wire  class_meta_rsp_fifo_io_in_bits_class_meta_field_type_19_is_repeated; // @[XQueue.scala 35:23]
  wire [4:0] class_meta_rsp_fifo_io_in_bits_class_meta_field_type_19_field_type; // @[XQueue.scala 35:23]
  wire [15:0] class_meta_rsp_fifo_io_in_bits_class_meta_field_type_19_sub_class_id; // @[XQueue.scala 35:23]
  wire  class_meta_rsp_fifo_io_in_bits_class_meta_field_type_20_is_repeated; // @[XQueue.scala 35:23]
  wire [4:0] class_meta_rsp_fifo_io_in_bits_class_meta_field_type_20_field_type; // @[XQueue.scala 35:23]
  wire [15:0] class_meta_rsp_fifo_io_in_bits_class_meta_field_type_20_sub_class_id; // @[XQueue.scala 35:23]
  wire  class_meta_rsp_fifo_io_in_bits_class_meta_field_type_21_is_repeated; // @[XQueue.scala 35:23]
  wire [4:0] class_meta_rsp_fifo_io_in_bits_class_meta_field_type_21_field_type; // @[XQueue.scala 35:23]
  wire [15:0] class_meta_rsp_fifo_io_in_bits_class_meta_field_type_21_sub_class_id; // @[XQueue.scala 35:23]
  wire  class_meta_rsp_fifo_io_in_bits_class_meta_field_type_22_is_repeated; // @[XQueue.scala 35:23]
  wire [4:0] class_meta_rsp_fifo_io_in_bits_class_meta_field_type_22_field_type; // @[XQueue.scala 35:23]
  wire [15:0] class_meta_rsp_fifo_io_in_bits_class_meta_field_type_22_sub_class_id; // @[XQueue.scala 35:23]
  wire  class_meta_rsp_fifo_io_in_bits_class_meta_field_type_23_is_repeated; // @[XQueue.scala 35:23]
  wire [4:0] class_meta_rsp_fifo_io_in_bits_class_meta_field_type_23_field_type; // @[XQueue.scala 35:23]
  wire [15:0] class_meta_rsp_fifo_io_in_bits_class_meta_field_type_23_sub_class_id; // @[XQueue.scala 35:23]
  wire  class_meta_rsp_fifo_io_in_bits_class_meta_field_type_24_is_repeated; // @[XQueue.scala 35:23]
  wire [4:0] class_meta_rsp_fifo_io_in_bits_class_meta_field_type_24_field_type; // @[XQueue.scala 35:23]
  wire [15:0] class_meta_rsp_fifo_io_in_bits_class_meta_field_type_24_sub_class_id; // @[XQueue.scala 35:23]
  wire  class_meta_rsp_fifo_io_in_bits_class_meta_field_type_25_is_repeated; // @[XQueue.scala 35:23]
  wire [4:0] class_meta_rsp_fifo_io_in_bits_class_meta_field_type_25_field_type; // @[XQueue.scala 35:23]
  wire [15:0] class_meta_rsp_fifo_io_in_bits_class_meta_field_type_25_sub_class_id; // @[XQueue.scala 35:23]
  wire  class_meta_rsp_fifo_io_in_bits_class_meta_field_type_26_is_repeated; // @[XQueue.scala 35:23]
  wire [4:0] class_meta_rsp_fifo_io_in_bits_class_meta_field_type_26_field_type; // @[XQueue.scala 35:23]
  wire [15:0] class_meta_rsp_fifo_io_in_bits_class_meta_field_type_26_sub_class_id; // @[XQueue.scala 35:23]
  wire  class_meta_rsp_fifo_io_in_bits_class_meta_field_type_27_is_repeated; // @[XQueue.scala 35:23]
  wire [4:0] class_meta_rsp_fifo_io_in_bits_class_meta_field_type_27_field_type; // @[XQueue.scala 35:23]
  wire [15:0] class_meta_rsp_fifo_io_in_bits_class_meta_field_type_27_sub_class_id; // @[XQueue.scala 35:23]
  wire  class_meta_rsp_fifo_io_in_bits_class_meta_field_type_28_is_repeated; // @[XQueue.scala 35:23]
  wire [4:0] class_meta_rsp_fifo_io_in_bits_class_meta_field_type_28_field_type; // @[XQueue.scala 35:23]
  wire [15:0] class_meta_rsp_fifo_io_in_bits_class_meta_field_type_28_sub_class_id; // @[XQueue.scala 35:23]
  wire  class_meta_rsp_fifo_io_in_bits_class_meta_field_type_29_is_repeated; // @[XQueue.scala 35:23]
  wire [4:0] class_meta_rsp_fifo_io_in_bits_class_meta_field_type_29_field_type; // @[XQueue.scala 35:23]
  wire [15:0] class_meta_rsp_fifo_io_in_bits_class_meta_field_type_29_sub_class_id; // @[XQueue.scala 35:23]
  wire  class_meta_rsp_fifo_io_in_bits_class_meta_field_type_30_is_repeated; // @[XQueue.scala 35:23]
  wire [4:0] class_meta_rsp_fifo_io_in_bits_class_meta_field_type_30_field_type; // @[XQueue.scala 35:23]
  wire [15:0] class_meta_rsp_fifo_io_in_bits_class_meta_field_type_30_sub_class_id; // @[XQueue.scala 35:23]
  wire  class_meta_rsp_fifo_io_in_bits_class_meta_field_type_31_is_repeated; // @[XQueue.scala 35:23]
  wire [4:0] class_meta_rsp_fifo_io_in_bits_class_meta_field_type_31_field_type; // @[XQueue.scala 35:23]
  wire [15:0] class_meta_rsp_fifo_io_in_bits_class_meta_field_type_31_sub_class_id; // @[XQueue.scala 35:23]
  wire  class_meta_rsp_fifo_io_in_bits_class_meta_field_type_32_is_repeated; // @[XQueue.scala 35:23]
  wire [4:0] class_meta_rsp_fifo_io_in_bits_class_meta_field_type_32_field_type; // @[XQueue.scala 35:23]
  wire [15:0] class_meta_rsp_fifo_io_in_bits_class_meta_field_type_32_sub_class_id; // @[XQueue.scala 35:23]
  wire  class_meta_rsp_fifo_io_out_ready; // @[XQueue.scala 35:23]
  wire  class_meta_rsp_fifo_io_out_valid; // @[XQueue.scala 35:23]
  wire [7:0] class_meta_rsp_fifo_io_out_bits_class_meta_max_field_num; // @[XQueue.scala 35:23]
  wire  class_meta_rsp_fifo_io_out_bits_class_meta_field_type_0_is_repeated; // @[XQueue.scala 35:23]
  wire [4:0] class_meta_rsp_fifo_io_out_bits_class_meta_field_type_0_field_type; // @[XQueue.scala 35:23]
  wire [15:0] class_meta_rsp_fifo_io_out_bits_class_meta_field_type_0_sub_class_id; // @[XQueue.scala 35:23]
  wire  class_meta_rsp_fifo_io_out_bits_class_meta_field_type_1_is_repeated; // @[XQueue.scala 35:23]
  wire [4:0] class_meta_rsp_fifo_io_out_bits_class_meta_field_type_1_field_type; // @[XQueue.scala 35:23]
  wire [15:0] class_meta_rsp_fifo_io_out_bits_class_meta_field_type_1_sub_class_id; // @[XQueue.scala 35:23]
  wire  class_meta_rsp_fifo_io_out_bits_class_meta_field_type_2_is_repeated; // @[XQueue.scala 35:23]
  wire [4:0] class_meta_rsp_fifo_io_out_bits_class_meta_field_type_2_field_type; // @[XQueue.scala 35:23]
  wire [15:0] class_meta_rsp_fifo_io_out_bits_class_meta_field_type_2_sub_class_id; // @[XQueue.scala 35:23]
  wire  class_meta_rsp_fifo_io_out_bits_class_meta_field_type_3_is_repeated; // @[XQueue.scala 35:23]
  wire [4:0] class_meta_rsp_fifo_io_out_bits_class_meta_field_type_3_field_type; // @[XQueue.scala 35:23]
  wire [15:0] class_meta_rsp_fifo_io_out_bits_class_meta_field_type_3_sub_class_id; // @[XQueue.scala 35:23]
  wire  class_meta_rsp_fifo_io_out_bits_class_meta_field_type_4_is_repeated; // @[XQueue.scala 35:23]
  wire [4:0] class_meta_rsp_fifo_io_out_bits_class_meta_field_type_4_field_type; // @[XQueue.scala 35:23]
  wire [15:0] class_meta_rsp_fifo_io_out_bits_class_meta_field_type_4_sub_class_id; // @[XQueue.scala 35:23]
  wire  class_meta_rsp_fifo_io_out_bits_class_meta_field_type_5_is_repeated; // @[XQueue.scala 35:23]
  wire [4:0] class_meta_rsp_fifo_io_out_bits_class_meta_field_type_5_field_type; // @[XQueue.scala 35:23]
  wire [15:0] class_meta_rsp_fifo_io_out_bits_class_meta_field_type_5_sub_class_id; // @[XQueue.scala 35:23]
  wire  class_meta_rsp_fifo_io_out_bits_class_meta_field_type_6_is_repeated; // @[XQueue.scala 35:23]
  wire [4:0] class_meta_rsp_fifo_io_out_bits_class_meta_field_type_6_field_type; // @[XQueue.scala 35:23]
  wire [15:0] class_meta_rsp_fifo_io_out_bits_class_meta_field_type_6_sub_class_id; // @[XQueue.scala 35:23]
  wire  class_meta_rsp_fifo_io_out_bits_class_meta_field_type_7_is_repeated; // @[XQueue.scala 35:23]
  wire [4:0] class_meta_rsp_fifo_io_out_bits_class_meta_field_type_7_field_type; // @[XQueue.scala 35:23]
  wire [15:0] class_meta_rsp_fifo_io_out_bits_class_meta_field_type_7_sub_class_id; // @[XQueue.scala 35:23]
  wire  class_meta_rsp_fifo_io_out_bits_class_meta_field_type_8_is_repeated; // @[XQueue.scala 35:23]
  wire [4:0] class_meta_rsp_fifo_io_out_bits_class_meta_field_type_8_field_type; // @[XQueue.scala 35:23]
  wire [15:0] class_meta_rsp_fifo_io_out_bits_class_meta_field_type_8_sub_class_id; // @[XQueue.scala 35:23]
  wire  class_meta_rsp_fifo_io_out_bits_class_meta_field_type_9_is_repeated; // @[XQueue.scala 35:23]
  wire [4:0] class_meta_rsp_fifo_io_out_bits_class_meta_field_type_9_field_type; // @[XQueue.scala 35:23]
  wire [15:0] class_meta_rsp_fifo_io_out_bits_class_meta_field_type_9_sub_class_id; // @[XQueue.scala 35:23]
  wire  class_meta_rsp_fifo_io_out_bits_class_meta_field_type_10_is_repeated; // @[XQueue.scala 35:23]
  wire [4:0] class_meta_rsp_fifo_io_out_bits_class_meta_field_type_10_field_type; // @[XQueue.scala 35:23]
  wire [15:0] class_meta_rsp_fifo_io_out_bits_class_meta_field_type_10_sub_class_id; // @[XQueue.scala 35:23]
  wire  class_meta_rsp_fifo_io_out_bits_class_meta_field_type_11_is_repeated; // @[XQueue.scala 35:23]
  wire [4:0] class_meta_rsp_fifo_io_out_bits_class_meta_field_type_11_field_type; // @[XQueue.scala 35:23]
  wire [15:0] class_meta_rsp_fifo_io_out_bits_class_meta_field_type_11_sub_class_id; // @[XQueue.scala 35:23]
  wire  class_meta_rsp_fifo_io_out_bits_class_meta_field_type_12_is_repeated; // @[XQueue.scala 35:23]
  wire [4:0] class_meta_rsp_fifo_io_out_bits_class_meta_field_type_12_field_type; // @[XQueue.scala 35:23]
  wire [15:0] class_meta_rsp_fifo_io_out_bits_class_meta_field_type_12_sub_class_id; // @[XQueue.scala 35:23]
  wire  class_meta_rsp_fifo_io_out_bits_class_meta_field_type_13_is_repeated; // @[XQueue.scala 35:23]
  wire [4:0] class_meta_rsp_fifo_io_out_bits_class_meta_field_type_13_field_type; // @[XQueue.scala 35:23]
  wire [15:0] class_meta_rsp_fifo_io_out_bits_class_meta_field_type_13_sub_class_id; // @[XQueue.scala 35:23]
  wire  class_meta_rsp_fifo_io_out_bits_class_meta_field_type_14_is_repeated; // @[XQueue.scala 35:23]
  wire [4:0] class_meta_rsp_fifo_io_out_bits_class_meta_field_type_14_field_type; // @[XQueue.scala 35:23]
  wire [15:0] class_meta_rsp_fifo_io_out_bits_class_meta_field_type_14_sub_class_id; // @[XQueue.scala 35:23]
  wire  class_meta_rsp_fifo_io_out_bits_class_meta_field_type_15_is_repeated; // @[XQueue.scala 35:23]
  wire [4:0] class_meta_rsp_fifo_io_out_bits_class_meta_field_type_15_field_type; // @[XQueue.scala 35:23]
  wire [15:0] class_meta_rsp_fifo_io_out_bits_class_meta_field_type_15_sub_class_id; // @[XQueue.scala 35:23]
  wire  class_meta_rsp_fifo_io_out_bits_class_meta_field_type_16_is_repeated; // @[XQueue.scala 35:23]
  wire [4:0] class_meta_rsp_fifo_io_out_bits_class_meta_field_type_16_field_type; // @[XQueue.scala 35:23]
  wire [15:0] class_meta_rsp_fifo_io_out_bits_class_meta_field_type_16_sub_class_id; // @[XQueue.scala 35:23]
  wire  class_meta_rsp_fifo_io_out_bits_class_meta_field_type_17_is_repeated; // @[XQueue.scala 35:23]
  wire [4:0] class_meta_rsp_fifo_io_out_bits_class_meta_field_type_17_field_type; // @[XQueue.scala 35:23]
  wire [15:0] class_meta_rsp_fifo_io_out_bits_class_meta_field_type_17_sub_class_id; // @[XQueue.scala 35:23]
  wire  class_meta_rsp_fifo_io_out_bits_class_meta_field_type_18_is_repeated; // @[XQueue.scala 35:23]
  wire [4:0] class_meta_rsp_fifo_io_out_bits_class_meta_field_type_18_field_type; // @[XQueue.scala 35:23]
  wire [15:0] class_meta_rsp_fifo_io_out_bits_class_meta_field_type_18_sub_class_id; // @[XQueue.scala 35:23]
  wire  class_meta_rsp_fifo_io_out_bits_class_meta_field_type_19_is_repeated; // @[XQueue.scala 35:23]
  wire [4:0] class_meta_rsp_fifo_io_out_bits_class_meta_field_type_19_field_type; // @[XQueue.scala 35:23]
  wire [15:0] class_meta_rsp_fifo_io_out_bits_class_meta_field_type_19_sub_class_id; // @[XQueue.scala 35:23]
  wire  class_meta_rsp_fifo_io_out_bits_class_meta_field_type_20_is_repeated; // @[XQueue.scala 35:23]
  wire [4:0] class_meta_rsp_fifo_io_out_bits_class_meta_field_type_20_field_type; // @[XQueue.scala 35:23]
  wire [15:0] class_meta_rsp_fifo_io_out_bits_class_meta_field_type_20_sub_class_id; // @[XQueue.scala 35:23]
  wire  class_meta_rsp_fifo_io_out_bits_class_meta_field_type_21_is_repeated; // @[XQueue.scala 35:23]
  wire [4:0] class_meta_rsp_fifo_io_out_bits_class_meta_field_type_21_field_type; // @[XQueue.scala 35:23]
  wire [15:0] class_meta_rsp_fifo_io_out_bits_class_meta_field_type_21_sub_class_id; // @[XQueue.scala 35:23]
  wire  class_meta_rsp_fifo_io_out_bits_class_meta_field_type_22_is_repeated; // @[XQueue.scala 35:23]
  wire [4:0] class_meta_rsp_fifo_io_out_bits_class_meta_field_type_22_field_type; // @[XQueue.scala 35:23]
  wire [15:0] class_meta_rsp_fifo_io_out_bits_class_meta_field_type_22_sub_class_id; // @[XQueue.scala 35:23]
  wire  class_meta_rsp_fifo_io_out_bits_class_meta_field_type_23_is_repeated; // @[XQueue.scala 35:23]
  wire [4:0] class_meta_rsp_fifo_io_out_bits_class_meta_field_type_23_field_type; // @[XQueue.scala 35:23]
  wire [15:0] class_meta_rsp_fifo_io_out_bits_class_meta_field_type_23_sub_class_id; // @[XQueue.scala 35:23]
  wire  class_meta_rsp_fifo_io_out_bits_class_meta_field_type_24_is_repeated; // @[XQueue.scala 35:23]
  wire [4:0] class_meta_rsp_fifo_io_out_bits_class_meta_field_type_24_field_type; // @[XQueue.scala 35:23]
  wire [15:0] class_meta_rsp_fifo_io_out_bits_class_meta_field_type_24_sub_class_id; // @[XQueue.scala 35:23]
  wire  class_meta_rsp_fifo_io_out_bits_class_meta_field_type_25_is_repeated; // @[XQueue.scala 35:23]
  wire [4:0] class_meta_rsp_fifo_io_out_bits_class_meta_field_type_25_field_type; // @[XQueue.scala 35:23]
  wire [15:0] class_meta_rsp_fifo_io_out_bits_class_meta_field_type_25_sub_class_id; // @[XQueue.scala 35:23]
  wire  class_meta_rsp_fifo_io_out_bits_class_meta_field_type_26_is_repeated; // @[XQueue.scala 35:23]
  wire [4:0] class_meta_rsp_fifo_io_out_bits_class_meta_field_type_26_field_type; // @[XQueue.scala 35:23]
  wire [15:0] class_meta_rsp_fifo_io_out_bits_class_meta_field_type_26_sub_class_id; // @[XQueue.scala 35:23]
  wire  class_meta_rsp_fifo_io_out_bits_class_meta_field_type_27_is_repeated; // @[XQueue.scala 35:23]
  wire [4:0] class_meta_rsp_fifo_io_out_bits_class_meta_field_type_27_field_type; // @[XQueue.scala 35:23]
  wire [15:0] class_meta_rsp_fifo_io_out_bits_class_meta_field_type_27_sub_class_id; // @[XQueue.scala 35:23]
  wire  class_meta_rsp_fifo_io_out_bits_class_meta_field_type_28_is_repeated; // @[XQueue.scala 35:23]
  wire [4:0] class_meta_rsp_fifo_io_out_bits_class_meta_field_type_28_field_type; // @[XQueue.scala 35:23]
  wire [15:0] class_meta_rsp_fifo_io_out_bits_class_meta_field_type_28_sub_class_id; // @[XQueue.scala 35:23]
  wire  class_meta_rsp_fifo_io_out_bits_class_meta_field_type_29_is_repeated; // @[XQueue.scala 35:23]
  wire [4:0] class_meta_rsp_fifo_io_out_bits_class_meta_field_type_29_field_type; // @[XQueue.scala 35:23]
  wire [15:0] class_meta_rsp_fifo_io_out_bits_class_meta_field_type_29_sub_class_id; // @[XQueue.scala 35:23]
  wire  class_meta_rsp_fifo_io_out_bits_class_meta_field_type_30_is_repeated; // @[XQueue.scala 35:23]
  wire [4:0] class_meta_rsp_fifo_io_out_bits_class_meta_field_type_30_field_type; // @[XQueue.scala 35:23]
  wire [15:0] class_meta_rsp_fifo_io_out_bits_class_meta_field_type_30_sub_class_id; // @[XQueue.scala 35:23]
  wire  class_meta_rsp_fifo_io_out_bits_class_meta_field_type_31_is_repeated; // @[XQueue.scala 35:23]
  wire [4:0] class_meta_rsp_fifo_io_out_bits_class_meta_field_type_31_field_type; // @[XQueue.scala 35:23]
  wire [15:0] class_meta_rsp_fifo_io_out_bits_class_meta_field_type_31_sub_class_id; // @[XQueue.scala 35:23]
  wire  class_meta_rsp_fifo_io_out_bits_class_meta_field_type_32_is_repeated; // @[XQueue.scala 35:23]
  wire [4:0] class_meta_rsp_fifo_io_out_bits_class_meta_field_type_32_field_type; // @[XQueue.scala 35:23]
  wire [15:0] class_meta_rsp_fifo_io_out_bits_class_meta_field_type_32_sub_class_id; // @[XQueue.scala 35:23]
  reg [31:0] counter; // @[Collector.scala 169:42]
  wire  _T = io_meta_in_ready & io_meta_in_valid; // @[Decoupled.scala 40:37]
  wire [31:0] _counter_T_1 = counter + 32'h1; // @[Collector.scala 171:51]
  reg [31:0] counter_1; // @[Collector.scala 169:42]
  wire  _T_1 = io_host_data_in_ready & io_host_data_in_valid; // @[Decoupled.scala 40:37]
  wire [31:0] _counter_T_3 = counter_1 + 32'h1; // @[Collector.scala 171:51]
  reg [31:0] counter_2; // @[Collector.scala 169:42]
  wire  _T_2 = io_host_data_cmd_ready & io_host_data_cmd_valid; // @[Decoupled.scala 40:37]
  wire [31:0] _counter_T_5 = counter_2 + 32'h1; // @[Collector.scala 171:51]
  reg [31:0] counter_3; // @[Collector.scala 169:42]
  wire [31:0] _counter_T_7 = counter_3 + 32'h1; // @[Collector.scala 171:51]
  reg  field_stack_0_field_type_0_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_0_field_type_0_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_0_field_type_0_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_0_field_type_1_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_0_field_type_1_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_0_field_type_1_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_0_field_type_2_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_0_field_type_2_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_0_field_type_2_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_0_field_type_3_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_0_field_type_3_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_0_field_type_3_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_0_field_type_4_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_0_field_type_4_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_0_field_type_4_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_0_field_type_5_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_0_field_type_5_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_0_field_type_5_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_0_field_type_6_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_0_field_type_6_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_0_field_type_6_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_0_field_type_7_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_0_field_type_7_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_0_field_type_7_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_0_field_type_8_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_0_field_type_8_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_0_field_type_8_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_0_field_type_9_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_0_field_type_9_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_0_field_type_9_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_0_field_type_10_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_0_field_type_10_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_0_field_type_10_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_0_field_type_11_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_0_field_type_11_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_0_field_type_11_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_0_field_type_12_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_0_field_type_12_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_0_field_type_12_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_0_field_type_13_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_0_field_type_13_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_0_field_type_13_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_0_field_type_14_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_0_field_type_14_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_0_field_type_14_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_0_field_type_15_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_0_field_type_15_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_0_field_type_15_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_0_field_type_16_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_0_field_type_16_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_0_field_type_16_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_0_field_type_17_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_0_field_type_17_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_0_field_type_17_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_0_field_type_18_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_0_field_type_18_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_0_field_type_18_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_0_field_type_19_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_0_field_type_19_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_0_field_type_19_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_0_field_type_20_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_0_field_type_20_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_0_field_type_20_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_0_field_type_21_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_0_field_type_21_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_0_field_type_21_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_0_field_type_22_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_0_field_type_22_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_0_field_type_22_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_0_field_type_23_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_0_field_type_23_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_0_field_type_23_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_0_field_type_24_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_0_field_type_24_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_0_field_type_24_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_0_field_type_25_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_0_field_type_25_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_0_field_type_25_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_0_field_type_26_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_0_field_type_26_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_0_field_type_26_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_0_field_type_27_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_0_field_type_27_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_0_field_type_27_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_0_field_type_28_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_0_field_type_28_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_0_field_type_28_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_0_field_type_29_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_0_field_type_29_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_0_field_type_29_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_0_field_type_30_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_0_field_type_30_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_0_field_type_30_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_0_field_type_31_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_0_field_type_31_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_0_field_type_31_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_0_field_type_32_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_0_field_type_32_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_0_field_type_32_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_1_field_type_0_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_1_field_type_0_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_1_field_type_0_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_1_field_type_1_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_1_field_type_1_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_1_field_type_1_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_1_field_type_2_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_1_field_type_2_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_1_field_type_2_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_1_field_type_3_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_1_field_type_3_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_1_field_type_3_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_1_field_type_4_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_1_field_type_4_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_1_field_type_4_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_1_field_type_5_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_1_field_type_5_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_1_field_type_5_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_1_field_type_6_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_1_field_type_6_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_1_field_type_6_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_1_field_type_7_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_1_field_type_7_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_1_field_type_7_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_1_field_type_8_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_1_field_type_8_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_1_field_type_8_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_1_field_type_9_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_1_field_type_9_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_1_field_type_9_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_1_field_type_10_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_1_field_type_10_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_1_field_type_10_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_1_field_type_11_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_1_field_type_11_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_1_field_type_11_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_1_field_type_12_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_1_field_type_12_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_1_field_type_12_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_1_field_type_13_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_1_field_type_13_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_1_field_type_13_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_1_field_type_14_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_1_field_type_14_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_1_field_type_14_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_1_field_type_15_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_1_field_type_15_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_1_field_type_15_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_1_field_type_16_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_1_field_type_16_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_1_field_type_16_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_1_field_type_17_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_1_field_type_17_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_1_field_type_17_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_1_field_type_18_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_1_field_type_18_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_1_field_type_18_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_1_field_type_19_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_1_field_type_19_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_1_field_type_19_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_1_field_type_20_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_1_field_type_20_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_1_field_type_20_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_1_field_type_21_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_1_field_type_21_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_1_field_type_21_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_1_field_type_22_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_1_field_type_22_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_1_field_type_22_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_1_field_type_23_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_1_field_type_23_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_1_field_type_23_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_1_field_type_24_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_1_field_type_24_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_1_field_type_24_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_1_field_type_25_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_1_field_type_25_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_1_field_type_25_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_1_field_type_26_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_1_field_type_26_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_1_field_type_26_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_1_field_type_27_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_1_field_type_27_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_1_field_type_27_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_1_field_type_28_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_1_field_type_28_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_1_field_type_28_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_1_field_type_29_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_1_field_type_29_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_1_field_type_29_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_1_field_type_30_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_1_field_type_30_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_1_field_type_30_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_1_field_type_31_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_1_field_type_31_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_1_field_type_31_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_1_field_type_32_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_1_field_type_32_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_1_field_type_32_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_2_field_type_0_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_2_field_type_0_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_2_field_type_0_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_2_field_type_1_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_2_field_type_1_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_2_field_type_1_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_2_field_type_2_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_2_field_type_2_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_2_field_type_2_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_2_field_type_3_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_2_field_type_3_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_2_field_type_3_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_2_field_type_4_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_2_field_type_4_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_2_field_type_4_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_2_field_type_5_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_2_field_type_5_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_2_field_type_5_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_2_field_type_6_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_2_field_type_6_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_2_field_type_6_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_2_field_type_7_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_2_field_type_7_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_2_field_type_7_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_2_field_type_8_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_2_field_type_8_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_2_field_type_8_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_2_field_type_9_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_2_field_type_9_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_2_field_type_9_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_2_field_type_10_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_2_field_type_10_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_2_field_type_10_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_2_field_type_11_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_2_field_type_11_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_2_field_type_11_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_2_field_type_12_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_2_field_type_12_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_2_field_type_12_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_2_field_type_13_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_2_field_type_13_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_2_field_type_13_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_2_field_type_14_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_2_field_type_14_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_2_field_type_14_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_2_field_type_15_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_2_field_type_15_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_2_field_type_15_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_2_field_type_16_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_2_field_type_16_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_2_field_type_16_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_2_field_type_17_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_2_field_type_17_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_2_field_type_17_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_2_field_type_18_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_2_field_type_18_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_2_field_type_18_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_2_field_type_19_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_2_field_type_19_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_2_field_type_19_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_2_field_type_20_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_2_field_type_20_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_2_field_type_20_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_2_field_type_21_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_2_field_type_21_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_2_field_type_21_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_2_field_type_22_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_2_field_type_22_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_2_field_type_22_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_2_field_type_23_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_2_field_type_23_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_2_field_type_23_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_2_field_type_24_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_2_field_type_24_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_2_field_type_24_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_2_field_type_25_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_2_field_type_25_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_2_field_type_25_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_2_field_type_26_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_2_field_type_26_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_2_field_type_26_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_2_field_type_27_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_2_field_type_27_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_2_field_type_27_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_2_field_type_28_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_2_field_type_28_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_2_field_type_28_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_2_field_type_29_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_2_field_type_29_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_2_field_type_29_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_2_field_type_30_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_2_field_type_30_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_2_field_type_30_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_2_field_type_31_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_2_field_type_31_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_2_field_type_31_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_2_field_type_32_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_2_field_type_32_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_2_field_type_32_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_3_field_type_0_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_3_field_type_0_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_3_field_type_0_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_3_field_type_1_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_3_field_type_1_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_3_field_type_1_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_3_field_type_2_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_3_field_type_2_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_3_field_type_2_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_3_field_type_3_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_3_field_type_3_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_3_field_type_3_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_3_field_type_4_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_3_field_type_4_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_3_field_type_4_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_3_field_type_5_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_3_field_type_5_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_3_field_type_5_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_3_field_type_6_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_3_field_type_6_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_3_field_type_6_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_3_field_type_7_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_3_field_type_7_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_3_field_type_7_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_3_field_type_8_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_3_field_type_8_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_3_field_type_8_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_3_field_type_9_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_3_field_type_9_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_3_field_type_9_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_3_field_type_10_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_3_field_type_10_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_3_field_type_10_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_3_field_type_11_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_3_field_type_11_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_3_field_type_11_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_3_field_type_12_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_3_field_type_12_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_3_field_type_12_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_3_field_type_13_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_3_field_type_13_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_3_field_type_13_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_3_field_type_14_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_3_field_type_14_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_3_field_type_14_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_3_field_type_15_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_3_field_type_15_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_3_field_type_15_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_3_field_type_16_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_3_field_type_16_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_3_field_type_16_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_3_field_type_17_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_3_field_type_17_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_3_field_type_17_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_3_field_type_18_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_3_field_type_18_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_3_field_type_18_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_3_field_type_19_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_3_field_type_19_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_3_field_type_19_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_3_field_type_20_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_3_field_type_20_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_3_field_type_20_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_3_field_type_21_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_3_field_type_21_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_3_field_type_21_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_3_field_type_22_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_3_field_type_22_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_3_field_type_22_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_3_field_type_23_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_3_field_type_23_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_3_field_type_23_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_3_field_type_24_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_3_field_type_24_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_3_field_type_24_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_3_field_type_25_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_3_field_type_25_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_3_field_type_25_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_3_field_type_26_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_3_field_type_26_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_3_field_type_26_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_3_field_type_27_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_3_field_type_27_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_3_field_type_27_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_3_field_type_28_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_3_field_type_28_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_3_field_type_28_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_3_field_type_29_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_3_field_type_29_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_3_field_type_29_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_3_field_type_30_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_3_field_type_30_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_3_field_type_30_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_3_field_type_31_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_3_field_type_31_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_3_field_type_31_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_3_field_type_32_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_3_field_type_32_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_3_field_type_32_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_4_field_type_0_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_4_field_type_0_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_4_field_type_0_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_4_field_type_1_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_4_field_type_1_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_4_field_type_1_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_4_field_type_2_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_4_field_type_2_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_4_field_type_2_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_4_field_type_3_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_4_field_type_3_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_4_field_type_3_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_4_field_type_4_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_4_field_type_4_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_4_field_type_4_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_4_field_type_5_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_4_field_type_5_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_4_field_type_5_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_4_field_type_6_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_4_field_type_6_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_4_field_type_6_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_4_field_type_7_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_4_field_type_7_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_4_field_type_7_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_4_field_type_8_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_4_field_type_8_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_4_field_type_8_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_4_field_type_9_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_4_field_type_9_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_4_field_type_9_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_4_field_type_10_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_4_field_type_10_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_4_field_type_10_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_4_field_type_11_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_4_field_type_11_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_4_field_type_11_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_4_field_type_12_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_4_field_type_12_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_4_field_type_12_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_4_field_type_13_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_4_field_type_13_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_4_field_type_13_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_4_field_type_14_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_4_field_type_14_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_4_field_type_14_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_4_field_type_15_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_4_field_type_15_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_4_field_type_15_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_4_field_type_16_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_4_field_type_16_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_4_field_type_16_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_4_field_type_17_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_4_field_type_17_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_4_field_type_17_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_4_field_type_18_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_4_field_type_18_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_4_field_type_18_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_4_field_type_19_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_4_field_type_19_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_4_field_type_19_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_4_field_type_20_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_4_field_type_20_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_4_field_type_20_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_4_field_type_21_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_4_field_type_21_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_4_field_type_21_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_4_field_type_22_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_4_field_type_22_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_4_field_type_22_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_4_field_type_23_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_4_field_type_23_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_4_field_type_23_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_4_field_type_24_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_4_field_type_24_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_4_field_type_24_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_4_field_type_25_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_4_field_type_25_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_4_field_type_25_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_4_field_type_26_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_4_field_type_26_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_4_field_type_26_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_4_field_type_27_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_4_field_type_27_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_4_field_type_27_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_4_field_type_28_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_4_field_type_28_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_4_field_type_28_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_4_field_type_29_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_4_field_type_29_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_4_field_type_29_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_4_field_type_30_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_4_field_type_30_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_4_field_type_30_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_4_field_type_31_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_4_field_type_31_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_4_field_type_31_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_4_field_type_32_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_4_field_type_32_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_4_field_type_32_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_5_field_type_0_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_5_field_type_0_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_5_field_type_0_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_5_field_type_1_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_5_field_type_1_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_5_field_type_1_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_5_field_type_2_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_5_field_type_2_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_5_field_type_2_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_5_field_type_3_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_5_field_type_3_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_5_field_type_3_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_5_field_type_4_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_5_field_type_4_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_5_field_type_4_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_5_field_type_5_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_5_field_type_5_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_5_field_type_5_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_5_field_type_6_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_5_field_type_6_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_5_field_type_6_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_5_field_type_7_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_5_field_type_7_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_5_field_type_7_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_5_field_type_8_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_5_field_type_8_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_5_field_type_8_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_5_field_type_9_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_5_field_type_9_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_5_field_type_9_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_5_field_type_10_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_5_field_type_10_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_5_field_type_10_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_5_field_type_11_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_5_field_type_11_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_5_field_type_11_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_5_field_type_12_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_5_field_type_12_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_5_field_type_12_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_5_field_type_13_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_5_field_type_13_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_5_field_type_13_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_5_field_type_14_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_5_field_type_14_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_5_field_type_14_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_5_field_type_15_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_5_field_type_15_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_5_field_type_15_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_5_field_type_16_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_5_field_type_16_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_5_field_type_16_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_5_field_type_17_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_5_field_type_17_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_5_field_type_17_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_5_field_type_18_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_5_field_type_18_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_5_field_type_18_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_5_field_type_19_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_5_field_type_19_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_5_field_type_19_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_5_field_type_20_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_5_field_type_20_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_5_field_type_20_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_5_field_type_21_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_5_field_type_21_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_5_field_type_21_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_5_field_type_22_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_5_field_type_22_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_5_field_type_22_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_5_field_type_23_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_5_field_type_23_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_5_field_type_23_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_5_field_type_24_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_5_field_type_24_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_5_field_type_24_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_5_field_type_25_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_5_field_type_25_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_5_field_type_25_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_5_field_type_26_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_5_field_type_26_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_5_field_type_26_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_5_field_type_27_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_5_field_type_27_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_5_field_type_27_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_5_field_type_28_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_5_field_type_28_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_5_field_type_28_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_5_field_type_29_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_5_field_type_29_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_5_field_type_29_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_5_field_type_30_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_5_field_type_30_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_5_field_type_30_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_5_field_type_31_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_5_field_type_31_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_5_field_type_31_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_5_field_type_32_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_5_field_type_32_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_5_field_type_32_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_6_field_type_0_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_6_field_type_0_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_6_field_type_0_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_6_field_type_1_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_6_field_type_1_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_6_field_type_1_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_6_field_type_2_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_6_field_type_2_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_6_field_type_2_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_6_field_type_3_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_6_field_type_3_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_6_field_type_3_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_6_field_type_4_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_6_field_type_4_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_6_field_type_4_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_6_field_type_5_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_6_field_type_5_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_6_field_type_5_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_6_field_type_6_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_6_field_type_6_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_6_field_type_6_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_6_field_type_7_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_6_field_type_7_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_6_field_type_7_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_6_field_type_8_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_6_field_type_8_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_6_field_type_8_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_6_field_type_9_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_6_field_type_9_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_6_field_type_9_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_6_field_type_10_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_6_field_type_10_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_6_field_type_10_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_6_field_type_11_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_6_field_type_11_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_6_field_type_11_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_6_field_type_12_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_6_field_type_12_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_6_field_type_12_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_6_field_type_13_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_6_field_type_13_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_6_field_type_13_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_6_field_type_14_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_6_field_type_14_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_6_field_type_14_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_6_field_type_15_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_6_field_type_15_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_6_field_type_15_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_6_field_type_16_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_6_field_type_16_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_6_field_type_16_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_6_field_type_17_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_6_field_type_17_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_6_field_type_17_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_6_field_type_18_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_6_field_type_18_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_6_field_type_18_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_6_field_type_19_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_6_field_type_19_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_6_field_type_19_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_6_field_type_20_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_6_field_type_20_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_6_field_type_20_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_6_field_type_21_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_6_field_type_21_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_6_field_type_21_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_6_field_type_22_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_6_field_type_22_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_6_field_type_22_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_6_field_type_23_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_6_field_type_23_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_6_field_type_23_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_6_field_type_24_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_6_field_type_24_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_6_field_type_24_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_6_field_type_25_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_6_field_type_25_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_6_field_type_25_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_6_field_type_26_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_6_field_type_26_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_6_field_type_26_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_6_field_type_27_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_6_field_type_27_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_6_field_type_27_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_6_field_type_28_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_6_field_type_28_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_6_field_type_28_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_6_field_type_29_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_6_field_type_29_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_6_field_type_29_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_6_field_type_30_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_6_field_type_30_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_6_field_type_30_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_6_field_type_31_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_6_field_type_31_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_6_field_type_31_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_6_field_type_32_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_6_field_type_32_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_6_field_type_32_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_7_field_type_0_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_7_field_type_0_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_7_field_type_0_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_7_field_type_1_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_7_field_type_1_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_7_field_type_1_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_7_field_type_2_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_7_field_type_2_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_7_field_type_2_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_7_field_type_3_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_7_field_type_3_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_7_field_type_3_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_7_field_type_4_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_7_field_type_4_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_7_field_type_4_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_7_field_type_5_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_7_field_type_5_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_7_field_type_5_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_7_field_type_6_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_7_field_type_6_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_7_field_type_6_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_7_field_type_7_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_7_field_type_7_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_7_field_type_7_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_7_field_type_8_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_7_field_type_8_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_7_field_type_8_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_7_field_type_9_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_7_field_type_9_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_7_field_type_9_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_7_field_type_10_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_7_field_type_10_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_7_field_type_10_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_7_field_type_11_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_7_field_type_11_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_7_field_type_11_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_7_field_type_12_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_7_field_type_12_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_7_field_type_12_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_7_field_type_13_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_7_field_type_13_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_7_field_type_13_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_7_field_type_14_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_7_field_type_14_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_7_field_type_14_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_7_field_type_15_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_7_field_type_15_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_7_field_type_15_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_7_field_type_16_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_7_field_type_16_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_7_field_type_16_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_7_field_type_17_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_7_field_type_17_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_7_field_type_17_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_7_field_type_18_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_7_field_type_18_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_7_field_type_18_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_7_field_type_19_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_7_field_type_19_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_7_field_type_19_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_7_field_type_20_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_7_field_type_20_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_7_field_type_20_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_7_field_type_21_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_7_field_type_21_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_7_field_type_21_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_7_field_type_22_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_7_field_type_22_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_7_field_type_22_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_7_field_type_23_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_7_field_type_23_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_7_field_type_23_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_7_field_type_24_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_7_field_type_24_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_7_field_type_24_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_7_field_type_25_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_7_field_type_25_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_7_field_type_25_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_7_field_type_26_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_7_field_type_26_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_7_field_type_26_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_7_field_type_27_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_7_field_type_27_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_7_field_type_27_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_7_field_type_28_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_7_field_type_28_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_7_field_type_28_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_7_field_type_29_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_7_field_type_29_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_7_field_type_29_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_7_field_type_30_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_7_field_type_30_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_7_field_type_30_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_7_field_type_31_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_7_field_type_31_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_7_field_type_31_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_7_field_type_32_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_7_field_type_32_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_7_field_type_32_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_8_field_type_0_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_8_field_type_0_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_8_field_type_0_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_8_field_type_1_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_8_field_type_1_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_8_field_type_1_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_8_field_type_2_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_8_field_type_2_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_8_field_type_2_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_8_field_type_3_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_8_field_type_3_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_8_field_type_3_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_8_field_type_4_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_8_field_type_4_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_8_field_type_4_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_8_field_type_5_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_8_field_type_5_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_8_field_type_5_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_8_field_type_6_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_8_field_type_6_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_8_field_type_6_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_8_field_type_7_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_8_field_type_7_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_8_field_type_7_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_8_field_type_8_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_8_field_type_8_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_8_field_type_8_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_8_field_type_9_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_8_field_type_9_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_8_field_type_9_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_8_field_type_10_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_8_field_type_10_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_8_field_type_10_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_8_field_type_11_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_8_field_type_11_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_8_field_type_11_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_8_field_type_12_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_8_field_type_12_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_8_field_type_12_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_8_field_type_13_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_8_field_type_13_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_8_field_type_13_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_8_field_type_14_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_8_field_type_14_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_8_field_type_14_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_8_field_type_15_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_8_field_type_15_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_8_field_type_15_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_8_field_type_16_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_8_field_type_16_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_8_field_type_16_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_8_field_type_17_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_8_field_type_17_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_8_field_type_17_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_8_field_type_18_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_8_field_type_18_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_8_field_type_18_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_8_field_type_19_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_8_field_type_19_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_8_field_type_19_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_8_field_type_20_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_8_field_type_20_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_8_field_type_20_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_8_field_type_21_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_8_field_type_21_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_8_field_type_21_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_8_field_type_22_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_8_field_type_22_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_8_field_type_22_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_8_field_type_23_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_8_field_type_23_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_8_field_type_23_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_8_field_type_24_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_8_field_type_24_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_8_field_type_24_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_8_field_type_25_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_8_field_type_25_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_8_field_type_25_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_8_field_type_26_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_8_field_type_26_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_8_field_type_26_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_8_field_type_27_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_8_field_type_27_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_8_field_type_27_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_8_field_type_28_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_8_field_type_28_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_8_field_type_28_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_8_field_type_29_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_8_field_type_29_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_8_field_type_29_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_8_field_type_30_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_8_field_type_30_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_8_field_type_30_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_8_field_type_31_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_8_field_type_31_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_8_field_type_31_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_8_field_type_32_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_8_field_type_32_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_8_field_type_32_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_9_field_type_0_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_9_field_type_0_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_9_field_type_0_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_9_field_type_1_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_9_field_type_1_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_9_field_type_1_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_9_field_type_2_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_9_field_type_2_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_9_field_type_2_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_9_field_type_3_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_9_field_type_3_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_9_field_type_3_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_9_field_type_4_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_9_field_type_4_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_9_field_type_4_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_9_field_type_5_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_9_field_type_5_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_9_field_type_5_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_9_field_type_6_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_9_field_type_6_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_9_field_type_6_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_9_field_type_7_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_9_field_type_7_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_9_field_type_7_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_9_field_type_8_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_9_field_type_8_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_9_field_type_8_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_9_field_type_9_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_9_field_type_9_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_9_field_type_9_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_9_field_type_10_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_9_field_type_10_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_9_field_type_10_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_9_field_type_11_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_9_field_type_11_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_9_field_type_11_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_9_field_type_12_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_9_field_type_12_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_9_field_type_12_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_9_field_type_13_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_9_field_type_13_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_9_field_type_13_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_9_field_type_14_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_9_field_type_14_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_9_field_type_14_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_9_field_type_15_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_9_field_type_15_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_9_field_type_15_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_9_field_type_16_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_9_field_type_16_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_9_field_type_16_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_9_field_type_17_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_9_field_type_17_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_9_field_type_17_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_9_field_type_18_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_9_field_type_18_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_9_field_type_18_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_9_field_type_19_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_9_field_type_19_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_9_field_type_19_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_9_field_type_20_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_9_field_type_20_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_9_field_type_20_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_9_field_type_21_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_9_field_type_21_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_9_field_type_21_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_9_field_type_22_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_9_field_type_22_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_9_field_type_22_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_9_field_type_23_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_9_field_type_23_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_9_field_type_23_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_9_field_type_24_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_9_field_type_24_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_9_field_type_24_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_9_field_type_25_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_9_field_type_25_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_9_field_type_25_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_9_field_type_26_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_9_field_type_26_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_9_field_type_26_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_9_field_type_27_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_9_field_type_27_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_9_field_type_27_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_9_field_type_28_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_9_field_type_28_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_9_field_type_28_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_9_field_type_29_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_9_field_type_29_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_9_field_type_29_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_9_field_type_30_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_9_field_type_30_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_9_field_type_30_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_9_field_type_31_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_9_field_type_31_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_9_field_type_31_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_9_field_type_32_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_9_field_type_32_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_9_field_type_32_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_10_field_type_0_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_10_field_type_0_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_10_field_type_0_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_10_field_type_1_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_10_field_type_1_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_10_field_type_1_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_10_field_type_2_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_10_field_type_2_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_10_field_type_2_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_10_field_type_3_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_10_field_type_3_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_10_field_type_3_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_10_field_type_4_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_10_field_type_4_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_10_field_type_4_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_10_field_type_5_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_10_field_type_5_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_10_field_type_5_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_10_field_type_6_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_10_field_type_6_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_10_field_type_6_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_10_field_type_7_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_10_field_type_7_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_10_field_type_7_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_10_field_type_8_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_10_field_type_8_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_10_field_type_8_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_10_field_type_9_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_10_field_type_9_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_10_field_type_9_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_10_field_type_10_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_10_field_type_10_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_10_field_type_10_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_10_field_type_11_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_10_field_type_11_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_10_field_type_11_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_10_field_type_12_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_10_field_type_12_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_10_field_type_12_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_10_field_type_13_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_10_field_type_13_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_10_field_type_13_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_10_field_type_14_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_10_field_type_14_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_10_field_type_14_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_10_field_type_15_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_10_field_type_15_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_10_field_type_15_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_10_field_type_16_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_10_field_type_16_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_10_field_type_16_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_10_field_type_17_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_10_field_type_17_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_10_field_type_17_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_10_field_type_18_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_10_field_type_18_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_10_field_type_18_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_10_field_type_19_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_10_field_type_19_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_10_field_type_19_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_10_field_type_20_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_10_field_type_20_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_10_field_type_20_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_10_field_type_21_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_10_field_type_21_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_10_field_type_21_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_10_field_type_22_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_10_field_type_22_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_10_field_type_22_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_10_field_type_23_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_10_field_type_23_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_10_field_type_23_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_10_field_type_24_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_10_field_type_24_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_10_field_type_24_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_10_field_type_25_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_10_field_type_25_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_10_field_type_25_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_10_field_type_26_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_10_field_type_26_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_10_field_type_26_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_10_field_type_27_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_10_field_type_27_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_10_field_type_27_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_10_field_type_28_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_10_field_type_28_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_10_field_type_28_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_10_field_type_29_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_10_field_type_29_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_10_field_type_29_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_10_field_type_30_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_10_field_type_30_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_10_field_type_30_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_10_field_type_31_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_10_field_type_31_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_10_field_type_31_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_10_field_type_32_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_10_field_type_32_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_10_field_type_32_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_11_field_type_0_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_11_field_type_0_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_11_field_type_0_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_11_field_type_1_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_11_field_type_1_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_11_field_type_1_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_11_field_type_2_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_11_field_type_2_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_11_field_type_2_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_11_field_type_3_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_11_field_type_3_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_11_field_type_3_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_11_field_type_4_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_11_field_type_4_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_11_field_type_4_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_11_field_type_5_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_11_field_type_5_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_11_field_type_5_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_11_field_type_6_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_11_field_type_6_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_11_field_type_6_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_11_field_type_7_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_11_field_type_7_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_11_field_type_7_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_11_field_type_8_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_11_field_type_8_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_11_field_type_8_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_11_field_type_9_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_11_field_type_9_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_11_field_type_9_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_11_field_type_10_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_11_field_type_10_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_11_field_type_10_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_11_field_type_11_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_11_field_type_11_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_11_field_type_11_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_11_field_type_12_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_11_field_type_12_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_11_field_type_12_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_11_field_type_13_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_11_field_type_13_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_11_field_type_13_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_11_field_type_14_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_11_field_type_14_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_11_field_type_14_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_11_field_type_15_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_11_field_type_15_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_11_field_type_15_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_11_field_type_16_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_11_field_type_16_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_11_field_type_16_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_11_field_type_17_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_11_field_type_17_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_11_field_type_17_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_11_field_type_18_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_11_field_type_18_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_11_field_type_18_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_11_field_type_19_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_11_field_type_19_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_11_field_type_19_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_11_field_type_20_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_11_field_type_20_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_11_field_type_20_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_11_field_type_21_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_11_field_type_21_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_11_field_type_21_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_11_field_type_22_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_11_field_type_22_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_11_field_type_22_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_11_field_type_23_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_11_field_type_23_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_11_field_type_23_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_11_field_type_24_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_11_field_type_24_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_11_field_type_24_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_11_field_type_25_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_11_field_type_25_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_11_field_type_25_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_11_field_type_26_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_11_field_type_26_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_11_field_type_26_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_11_field_type_27_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_11_field_type_27_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_11_field_type_27_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_11_field_type_28_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_11_field_type_28_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_11_field_type_28_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_11_field_type_29_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_11_field_type_29_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_11_field_type_29_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_11_field_type_30_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_11_field_type_30_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_11_field_type_30_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_11_field_type_31_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_11_field_type_31_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_11_field_type_31_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_11_field_type_32_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_11_field_type_32_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_11_field_type_32_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_12_field_type_0_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_12_field_type_0_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_12_field_type_0_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_12_field_type_1_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_12_field_type_1_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_12_field_type_1_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_12_field_type_2_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_12_field_type_2_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_12_field_type_2_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_12_field_type_3_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_12_field_type_3_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_12_field_type_3_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_12_field_type_4_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_12_field_type_4_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_12_field_type_4_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_12_field_type_5_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_12_field_type_5_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_12_field_type_5_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_12_field_type_6_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_12_field_type_6_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_12_field_type_6_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_12_field_type_7_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_12_field_type_7_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_12_field_type_7_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_12_field_type_8_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_12_field_type_8_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_12_field_type_8_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_12_field_type_9_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_12_field_type_9_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_12_field_type_9_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_12_field_type_10_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_12_field_type_10_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_12_field_type_10_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_12_field_type_11_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_12_field_type_11_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_12_field_type_11_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_12_field_type_12_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_12_field_type_12_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_12_field_type_12_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_12_field_type_13_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_12_field_type_13_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_12_field_type_13_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_12_field_type_14_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_12_field_type_14_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_12_field_type_14_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_12_field_type_15_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_12_field_type_15_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_12_field_type_15_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_12_field_type_16_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_12_field_type_16_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_12_field_type_16_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_12_field_type_17_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_12_field_type_17_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_12_field_type_17_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_12_field_type_18_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_12_field_type_18_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_12_field_type_18_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_12_field_type_19_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_12_field_type_19_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_12_field_type_19_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_12_field_type_20_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_12_field_type_20_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_12_field_type_20_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_12_field_type_21_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_12_field_type_21_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_12_field_type_21_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_12_field_type_22_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_12_field_type_22_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_12_field_type_22_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_12_field_type_23_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_12_field_type_23_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_12_field_type_23_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_12_field_type_24_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_12_field_type_24_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_12_field_type_24_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_12_field_type_25_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_12_field_type_25_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_12_field_type_25_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_12_field_type_26_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_12_field_type_26_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_12_field_type_26_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_12_field_type_27_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_12_field_type_27_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_12_field_type_27_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_12_field_type_28_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_12_field_type_28_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_12_field_type_28_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_12_field_type_29_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_12_field_type_29_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_12_field_type_29_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_12_field_type_30_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_12_field_type_30_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_12_field_type_30_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_12_field_type_31_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_12_field_type_31_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_12_field_type_31_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_12_field_type_32_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_12_field_type_32_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_12_field_type_32_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_13_field_type_0_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_13_field_type_0_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_13_field_type_0_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_13_field_type_1_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_13_field_type_1_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_13_field_type_1_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_13_field_type_2_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_13_field_type_2_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_13_field_type_2_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_13_field_type_3_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_13_field_type_3_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_13_field_type_3_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_13_field_type_4_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_13_field_type_4_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_13_field_type_4_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_13_field_type_5_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_13_field_type_5_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_13_field_type_5_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_13_field_type_6_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_13_field_type_6_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_13_field_type_6_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_13_field_type_7_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_13_field_type_7_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_13_field_type_7_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_13_field_type_8_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_13_field_type_8_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_13_field_type_8_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_13_field_type_9_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_13_field_type_9_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_13_field_type_9_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_13_field_type_10_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_13_field_type_10_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_13_field_type_10_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_13_field_type_11_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_13_field_type_11_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_13_field_type_11_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_13_field_type_12_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_13_field_type_12_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_13_field_type_12_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_13_field_type_13_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_13_field_type_13_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_13_field_type_13_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_13_field_type_14_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_13_field_type_14_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_13_field_type_14_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_13_field_type_15_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_13_field_type_15_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_13_field_type_15_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_13_field_type_16_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_13_field_type_16_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_13_field_type_16_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_13_field_type_17_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_13_field_type_17_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_13_field_type_17_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_13_field_type_18_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_13_field_type_18_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_13_field_type_18_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_13_field_type_19_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_13_field_type_19_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_13_field_type_19_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_13_field_type_20_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_13_field_type_20_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_13_field_type_20_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_13_field_type_21_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_13_field_type_21_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_13_field_type_21_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_13_field_type_22_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_13_field_type_22_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_13_field_type_22_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_13_field_type_23_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_13_field_type_23_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_13_field_type_23_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_13_field_type_24_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_13_field_type_24_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_13_field_type_24_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_13_field_type_25_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_13_field_type_25_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_13_field_type_25_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_13_field_type_26_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_13_field_type_26_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_13_field_type_26_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_13_field_type_27_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_13_field_type_27_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_13_field_type_27_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_13_field_type_28_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_13_field_type_28_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_13_field_type_28_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_13_field_type_29_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_13_field_type_29_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_13_field_type_29_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_13_field_type_30_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_13_field_type_30_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_13_field_type_30_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_13_field_type_31_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_13_field_type_31_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_13_field_type_31_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_13_field_type_32_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_13_field_type_32_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_13_field_type_32_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_14_field_type_0_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_14_field_type_0_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_14_field_type_0_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_14_field_type_1_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_14_field_type_1_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_14_field_type_1_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_14_field_type_2_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_14_field_type_2_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_14_field_type_2_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_14_field_type_3_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_14_field_type_3_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_14_field_type_3_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_14_field_type_4_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_14_field_type_4_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_14_field_type_4_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_14_field_type_5_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_14_field_type_5_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_14_field_type_5_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_14_field_type_6_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_14_field_type_6_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_14_field_type_6_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_14_field_type_7_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_14_field_type_7_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_14_field_type_7_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_14_field_type_8_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_14_field_type_8_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_14_field_type_8_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_14_field_type_9_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_14_field_type_9_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_14_field_type_9_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_14_field_type_10_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_14_field_type_10_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_14_field_type_10_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_14_field_type_11_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_14_field_type_11_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_14_field_type_11_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_14_field_type_12_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_14_field_type_12_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_14_field_type_12_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_14_field_type_13_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_14_field_type_13_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_14_field_type_13_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_14_field_type_14_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_14_field_type_14_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_14_field_type_14_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_14_field_type_15_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_14_field_type_15_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_14_field_type_15_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_14_field_type_16_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_14_field_type_16_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_14_field_type_16_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_14_field_type_17_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_14_field_type_17_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_14_field_type_17_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_14_field_type_18_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_14_field_type_18_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_14_field_type_18_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_14_field_type_19_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_14_field_type_19_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_14_field_type_19_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_14_field_type_20_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_14_field_type_20_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_14_field_type_20_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_14_field_type_21_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_14_field_type_21_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_14_field_type_21_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_14_field_type_22_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_14_field_type_22_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_14_field_type_22_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_14_field_type_23_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_14_field_type_23_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_14_field_type_23_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_14_field_type_24_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_14_field_type_24_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_14_field_type_24_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_14_field_type_25_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_14_field_type_25_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_14_field_type_25_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_14_field_type_26_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_14_field_type_26_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_14_field_type_26_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_14_field_type_27_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_14_field_type_27_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_14_field_type_27_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_14_field_type_28_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_14_field_type_28_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_14_field_type_28_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_14_field_type_29_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_14_field_type_29_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_14_field_type_29_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_14_field_type_30_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_14_field_type_30_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_14_field_type_30_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_14_field_type_31_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_14_field_type_31_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_14_field_type_31_sub_class_id; // @[Serializerhw.scala 68:30]
  reg  field_stack_14_field_type_32_is_repeated; // @[Serializerhw.scala 68:30]
  reg [4:0] field_stack_14_field_type_32_field_type; // @[Serializerhw.scala 68:30]
  reg [15:0] field_stack_14_field_type_32_sub_class_id; // @[Serializerhw.scala 68:30]
  reg [5:0] field_num_0; // @[Serializerhw.scala 70:28]
  reg [5:0] field_num_1; // @[Serializerhw.scala 70:28]
  reg [5:0] field_num_2; // @[Serializerhw.scala 70:28]
  reg [5:0] field_num_3; // @[Serializerhw.scala 70:28]
  reg [5:0] field_num_4; // @[Serializerhw.scala 70:28]
  reg [5:0] field_num_5; // @[Serializerhw.scala 70:28]
  reg [5:0] field_num_6; // @[Serializerhw.scala 70:28]
  reg [5:0] field_num_7; // @[Serializerhw.scala 70:28]
  reg [5:0] field_num_8; // @[Serializerhw.scala 70:28]
  reg [5:0] field_num_9; // @[Serializerhw.scala 70:28]
  reg [5:0] field_num_10; // @[Serializerhw.scala 70:28]
  reg [5:0] field_num_11; // @[Serializerhw.scala 70:28]
  reg [5:0] field_num_12; // @[Serializerhw.scala 70:28]
  reg [5:0] field_num_13; // @[Serializerhw.scala 70:28]
  reg [5:0] field_num_14; // @[Serializerhw.scala 70:28]
  reg [5:0] field_num_15; // @[Serializerhw.scala 70:28]
  reg [63:0] host_base_addr; // @[Serializerhw.scala 72:33]
  reg [5:0] current_field_num; // @[Serializerhw.scala 73:36]
  reg  c_sub_metadata_is_repeated; // @[Serializerhw.scala 74:33]
  reg [4:0] c_sub_metadata_field_type; // @[Serializerhw.scala 74:33]
  reg [15:0] c_sub_metadata_sub_class_id; // @[Serializerhw.scala 74:33]
  reg [7:0] repeat_num; // @[Serializerhw.scala 75:29]
  reg [3:0] stack_num; // @[Serializerhw.scala 76:30]
  reg [31:0] current_field_length; // @[Serializerhw.scala 83:38]
  reg [4:0] state; // @[Serializerhw.scala 86:46]
  wire  _T_4 = 5'h6 == state; // @[Conditional.scala 37:30]
  wire  _T_5 = meta_in_fifo_io_out_ready & meta_in_fifo_io_out_valid; // @[Decoupled.scala 40:37]
  wire [9:0] _GEN_12 = _T_5 ? meta_in_fifo_io_out_bits_class_id : 10'h0; // @[Serializerhw.scala 102:45 Serializerhw.scala 106:50 Util.scala 13:25]
  wire  _T_6 = 5'h11 == state; // @[Conditional.scala 37:30]
  wire  _T_7 = class_meta_rsp_fifo_io_out_ready & class_meta_rsp_fifo_io_out_valid; // @[Decoupled.scala 40:37]
  wire [15:0] _field_stack_stack_num_field_type_0_sub_class_id =
    class_meta_rsp_fifo_io_out_bits_class_meta_field_type_0_sub_class_id; // @[Serializerhw.scala 114:45 Serializerhw.scala 114:45]
  wire [4:0] _field_stack_stack_num_field_type_0_field_type =
    class_meta_rsp_fifo_io_out_bits_class_meta_field_type_0_field_type; // @[Serializerhw.scala 114:45 Serializerhw.scala 114:45]
  wire [15:0] _field_stack_stack_num_field_type_1_sub_class_id =
    class_meta_rsp_fifo_io_out_bits_class_meta_field_type_1_sub_class_id; // @[Serializerhw.scala 114:45 Serializerhw.scala 114:45]
  wire [4:0] _field_stack_stack_num_field_type_1_field_type =
    class_meta_rsp_fifo_io_out_bits_class_meta_field_type_1_field_type; // @[Serializerhw.scala 114:45 Serializerhw.scala 114:45]
  wire [15:0] _field_stack_stack_num_field_type_2_sub_class_id =
    class_meta_rsp_fifo_io_out_bits_class_meta_field_type_2_sub_class_id; // @[Serializerhw.scala 114:45 Serializerhw.scala 114:45]
  wire [4:0] _field_stack_stack_num_field_type_2_field_type =
    class_meta_rsp_fifo_io_out_bits_class_meta_field_type_2_field_type; // @[Serializerhw.scala 114:45 Serializerhw.scala 114:45]
  wire [15:0] _field_stack_stack_num_field_type_3_sub_class_id =
    class_meta_rsp_fifo_io_out_bits_class_meta_field_type_3_sub_class_id; // @[Serializerhw.scala 114:45 Serializerhw.scala 114:45]
  wire [4:0] _field_stack_stack_num_field_type_3_field_type =
    class_meta_rsp_fifo_io_out_bits_class_meta_field_type_3_field_type; // @[Serializerhw.scala 114:45 Serializerhw.scala 114:45]
  wire [15:0] _field_stack_stack_num_field_type_4_sub_class_id =
    class_meta_rsp_fifo_io_out_bits_class_meta_field_type_4_sub_class_id; // @[Serializerhw.scala 114:45 Serializerhw.scala 114:45]
  wire [4:0] _field_stack_stack_num_field_type_4_field_type =
    class_meta_rsp_fifo_io_out_bits_class_meta_field_type_4_field_type; // @[Serializerhw.scala 114:45 Serializerhw.scala 114:45]
  wire [15:0] _field_stack_stack_num_field_type_5_sub_class_id =
    class_meta_rsp_fifo_io_out_bits_class_meta_field_type_5_sub_class_id; // @[Serializerhw.scala 114:45 Serializerhw.scala 114:45]
  wire [4:0] _field_stack_stack_num_field_type_5_field_type =
    class_meta_rsp_fifo_io_out_bits_class_meta_field_type_5_field_type; // @[Serializerhw.scala 114:45 Serializerhw.scala 114:45]
  wire [15:0] _field_stack_stack_num_field_type_6_sub_class_id =
    class_meta_rsp_fifo_io_out_bits_class_meta_field_type_6_sub_class_id; // @[Serializerhw.scala 114:45 Serializerhw.scala 114:45]
  wire [4:0] _field_stack_stack_num_field_type_6_field_type =
    class_meta_rsp_fifo_io_out_bits_class_meta_field_type_6_field_type; // @[Serializerhw.scala 114:45 Serializerhw.scala 114:45]
  wire [15:0] _field_stack_stack_num_field_type_7_sub_class_id =
    class_meta_rsp_fifo_io_out_bits_class_meta_field_type_7_sub_class_id; // @[Serializerhw.scala 114:45 Serializerhw.scala 114:45]
  wire [4:0] _field_stack_stack_num_field_type_7_field_type =
    class_meta_rsp_fifo_io_out_bits_class_meta_field_type_7_field_type; // @[Serializerhw.scala 114:45 Serializerhw.scala 114:45]
  wire [15:0] _field_stack_stack_num_field_type_8_sub_class_id =
    class_meta_rsp_fifo_io_out_bits_class_meta_field_type_8_sub_class_id; // @[Serializerhw.scala 114:45 Serializerhw.scala 114:45]
  wire [4:0] _field_stack_stack_num_field_type_8_field_type =
    class_meta_rsp_fifo_io_out_bits_class_meta_field_type_8_field_type; // @[Serializerhw.scala 114:45 Serializerhw.scala 114:45]
  wire [15:0] _field_stack_stack_num_field_type_9_sub_class_id =
    class_meta_rsp_fifo_io_out_bits_class_meta_field_type_9_sub_class_id; // @[Serializerhw.scala 114:45 Serializerhw.scala 114:45]
  wire [4:0] _field_stack_stack_num_field_type_9_field_type =
    class_meta_rsp_fifo_io_out_bits_class_meta_field_type_9_field_type; // @[Serializerhw.scala 114:45 Serializerhw.scala 114:45]
  wire [15:0] _field_stack_stack_num_field_type_10_sub_class_id =
    class_meta_rsp_fifo_io_out_bits_class_meta_field_type_10_sub_class_id; // @[Serializerhw.scala 114:45 Serializerhw.scala 114:45]
  wire [4:0] _field_stack_stack_num_field_type_10_field_type =
    class_meta_rsp_fifo_io_out_bits_class_meta_field_type_10_field_type; // @[Serializerhw.scala 114:45 Serializerhw.scala 114:45]
  wire [15:0] _field_stack_stack_num_field_type_11_sub_class_id =
    class_meta_rsp_fifo_io_out_bits_class_meta_field_type_11_sub_class_id; // @[Serializerhw.scala 114:45 Serializerhw.scala 114:45]
  wire [4:0] _field_stack_stack_num_field_type_11_field_type =
    class_meta_rsp_fifo_io_out_bits_class_meta_field_type_11_field_type; // @[Serializerhw.scala 114:45 Serializerhw.scala 114:45]
  wire [15:0] _field_stack_stack_num_field_type_12_sub_class_id =
    class_meta_rsp_fifo_io_out_bits_class_meta_field_type_12_sub_class_id; // @[Serializerhw.scala 114:45 Serializerhw.scala 114:45]
  wire [4:0] _field_stack_stack_num_field_type_12_field_type =
    class_meta_rsp_fifo_io_out_bits_class_meta_field_type_12_field_type; // @[Serializerhw.scala 114:45 Serializerhw.scala 114:45]
  wire [15:0] _field_stack_stack_num_field_type_13_sub_class_id =
    class_meta_rsp_fifo_io_out_bits_class_meta_field_type_13_sub_class_id; // @[Serializerhw.scala 114:45 Serializerhw.scala 114:45]
  wire [4:0] _field_stack_stack_num_field_type_13_field_type =
    class_meta_rsp_fifo_io_out_bits_class_meta_field_type_13_field_type; // @[Serializerhw.scala 114:45 Serializerhw.scala 114:45]
  wire [15:0] _field_stack_stack_num_field_type_14_sub_class_id =
    class_meta_rsp_fifo_io_out_bits_class_meta_field_type_14_sub_class_id; // @[Serializerhw.scala 114:45 Serializerhw.scala 114:45]
  wire [4:0] _field_stack_stack_num_field_type_14_field_type =
    class_meta_rsp_fifo_io_out_bits_class_meta_field_type_14_field_type; // @[Serializerhw.scala 114:45 Serializerhw.scala 114:45]
  wire [15:0] _field_stack_stack_num_field_type_15_sub_class_id =
    class_meta_rsp_fifo_io_out_bits_class_meta_field_type_15_sub_class_id; // @[Serializerhw.scala 114:45 Serializerhw.scala 114:45]
  wire [4:0] _field_stack_stack_num_field_type_15_field_type =
    class_meta_rsp_fifo_io_out_bits_class_meta_field_type_15_field_type; // @[Serializerhw.scala 114:45 Serializerhw.scala 114:45]
  wire [15:0] _field_stack_stack_num_field_type_16_sub_class_id =
    class_meta_rsp_fifo_io_out_bits_class_meta_field_type_16_sub_class_id; // @[Serializerhw.scala 114:45 Serializerhw.scala 114:45]
  wire [4:0] _field_stack_stack_num_field_type_16_field_type =
    class_meta_rsp_fifo_io_out_bits_class_meta_field_type_16_field_type; // @[Serializerhw.scala 114:45 Serializerhw.scala 114:45]
  wire [15:0] _field_stack_stack_num_field_type_17_sub_class_id =
    class_meta_rsp_fifo_io_out_bits_class_meta_field_type_17_sub_class_id; // @[Serializerhw.scala 114:45 Serializerhw.scala 114:45]
  wire [4:0] _field_stack_stack_num_field_type_17_field_type =
    class_meta_rsp_fifo_io_out_bits_class_meta_field_type_17_field_type; // @[Serializerhw.scala 114:45 Serializerhw.scala 114:45]
  wire [15:0] _field_stack_stack_num_field_type_18_sub_class_id =
    class_meta_rsp_fifo_io_out_bits_class_meta_field_type_18_sub_class_id; // @[Serializerhw.scala 114:45 Serializerhw.scala 114:45]
  wire [4:0] _field_stack_stack_num_field_type_18_field_type =
    class_meta_rsp_fifo_io_out_bits_class_meta_field_type_18_field_type; // @[Serializerhw.scala 114:45 Serializerhw.scala 114:45]
  wire [15:0] _field_stack_stack_num_field_type_19_sub_class_id =
    class_meta_rsp_fifo_io_out_bits_class_meta_field_type_19_sub_class_id; // @[Serializerhw.scala 114:45 Serializerhw.scala 114:45]
  wire [4:0] _field_stack_stack_num_field_type_19_field_type =
    class_meta_rsp_fifo_io_out_bits_class_meta_field_type_19_field_type; // @[Serializerhw.scala 114:45 Serializerhw.scala 114:45]
  wire [15:0] _field_stack_stack_num_field_type_20_sub_class_id =
    class_meta_rsp_fifo_io_out_bits_class_meta_field_type_20_sub_class_id; // @[Serializerhw.scala 114:45 Serializerhw.scala 114:45]
  wire [4:0] _field_stack_stack_num_field_type_20_field_type =
    class_meta_rsp_fifo_io_out_bits_class_meta_field_type_20_field_type; // @[Serializerhw.scala 114:45 Serializerhw.scala 114:45]
  wire [15:0] _field_stack_stack_num_field_type_21_sub_class_id =
    class_meta_rsp_fifo_io_out_bits_class_meta_field_type_21_sub_class_id; // @[Serializerhw.scala 114:45 Serializerhw.scala 114:45]
  wire [4:0] _field_stack_stack_num_field_type_21_field_type =
    class_meta_rsp_fifo_io_out_bits_class_meta_field_type_21_field_type; // @[Serializerhw.scala 114:45 Serializerhw.scala 114:45]
  wire [15:0] _field_stack_stack_num_field_type_22_sub_class_id =
    class_meta_rsp_fifo_io_out_bits_class_meta_field_type_22_sub_class_id; // @[Serializerhw.scala 114:45 Serializerhw.scala 114:45]
  wire [4:0] _field_stack_stack_num_field_type_22_field_type =
    class_meta_rsp_fifo_io_out_bits_class_meta_field_type_22_field_type; // @[Serializerhw.scala 114:45 Serializerhw.scala 114:45]
  wire [15:0] _field_stack_stack_num_field_type_23_sub_class_id =
    class_meta_rsp_fifo_io_out_bits_class_meta_field_type_23_sub_class_id; // @[Serializerhw.scala 114:45 Serializerhw.scala 114:45]
  wire [4:0] _field_stack_stack_num_field_type_23_field_type =
    class_meta_rsp_fifo_io_out_bits_class_meta_field_type_23_field_type; // @[Serializerhw.scala 114:45 Serializerhw.scala 114:45]
  wire [15:0] _field_stack_stack_num_field_type_24_sub_class_id =
    class_meta_rsp_fifo_io_out_bits_class_meta_field_type_24_sub_class_id; // @[Serializerhw.scala 114:45 Serializerhw.scala 114:45]
  wire [4:0] _field_stack_stack_num_field_type_24_field_type =
    class_meta_rsp_fifo_io_out_bits_class_meta_field_type_24_field_type; // @[Serializerhw.scala 114:45 Serializerhw.scala 114:45]
  wire [15:0] _field_stack_stack_num_field_type_25_sub_class_id =
    class_meta_rsp_fifo_io_out_bits_class_meta_field_type_25_sub_class_id; // @[Serializerhw.scala 114:45 Serializerhw.scala 114:45]
  wire [4:0] _field_stack_stack_num_field_type_25_field_type =
    class_meta_rsp_fifo_io_out_bits_class_meta_field_type_25_field_type; // @[Serializerhw.scala 114:45 Serializerhw.scala 114:45]
  wire [15:0] _field_stack_stack_num_field_type_26_sub_class_id =
    class_meta_rsp_fifo_io_out_bits_class_meta_field_type_26_sub_class_id; // @[Serializerhw.scala 114:45 Serializerhw.scala 114:45]
  wire [4:0] _field_stack_stack_num_field_type_26_field_type =
    class_meta_rsp_fifo_io_out_bits_class_meta_field_type_26_field_type; // @[Serializerhw.scala 114:45 Serializerhw.scala 114:45]
  wire [15:0] _field_stack_stack_num_field_type_27_sub_class_id =
    class_meta_rsp_fifo_io_out_bits_class_meta_field_type_27_sub_class_id; // @[Serializerhw.scala 114:45 Serializerhw.scala 114:45]
  wire [4:0] _field_stack_stack_num_field_type_27_field_type =
    class_meta_rsp_fifo_io_out_bits_class_meta_field_type_27_field_type; // @[Serializerhw.scala 114:45 Serializerhw.scala 114:45]
  wire [15:0] _field_stack_stack_num_field_type_28_sub_class_id =
    class_meta_rsp_fifo_io_out_bits_class_meta_field_type_28_sub_class_id; // @[Serializerhw.scala 114:45 Serializerhw.scala 114:45]
  wire [4:0] _field_stack_stack_num_field_type_28_field_type =
    class_meta_rsp_fifo_io_out_bits_class_meta_field_type_28_field_type; // @[Serializerhw.scala 114:45 Serializerhw.scala 114:45]
  wire [15:0] _field_stack_stack_num_field_type_29_sub_class_id =
    class_meta_rsp_fifo_io_out_bits_class_meta_field_type_29_sub_class_id; // @[Serializerhw.scala 114:45 Serializerhw.scala 114:45]
  wire [4:0] _field_stack_stack_num_field_type_29_field_type =
    class_meta_rsp_fifo_io_out_bits_class_meta_field_type_29_field_type; // @[Serializerhw.scala 114:45 Serializerhw.scala 114:45]
  wire [15:0] _field_stack_stack_num_field_type_30_sub_class_id =
    class_meta_rsp_fifo_io_out_bits_class_meta_field_type_30_sub_class_id; // @[Serializerhw.scala 114:45 Serializerhw.scala 114:45]
  wire [4:0] _field_stack_stack_num_field_type_30_field_type =
    class_meta_rsp_fifo_io_out_bits_class_meta_field_type_30_field_type; // @[Serializerhw.scala 114:45 Serializerhw.scala 114:45]
  wire [15:0] _field_stack_stack_num_field_type_31_sub_class_id =
    class_meta_rsp_fifo_io_out_bits_class_meta_field_type_31_sub_class_id; // @[Serializerhw.scala 114:45 Serializerhw.scala 114:45]
  wire [4:0] _field_stack_stack_num_field_type_31_field_type =
    class_meta_rsp_fifo_io_out_bits_class_meta_field_type_31_field_type; // @[Serializerhw.scala 114:45 Serializerhw.scala 114:45]
  wire [15:0] _field_stack_stack_num_field_type_32_sub_class_id =
    class_meta_rsp_fifo_io_out_bits_class_meta_field_type_32_sub_class_id; // @[Serializerhw.scala 114:45 Serializerhw.scala 114:45]
  wire [4:0] _field_stack_stack_num_field_type_32_field_type =
    class_meta_rsp_fifo_io_out_bits_class_meta_field_type_32_field_type; // @[Serializerhw.scala 114:45 Serializerhw.scala 114:45]
  wire [5:0] _GEN_2026 = 4'h0 == stack_num ? class_meta_rsp_fifo_io_out_bits_class_meta_max_field_num[5:0] : field_num_0
    ; // @[Serializerhw.scala 115:45 Serializerhw.scala 115:45 Serializerhw.scala 70:28]
  wire [5:0] _GEN_2027 = 4'h1 == stack_num ? class_meta_rsp_fifo_io_out_bits_class_meta_max_field_num[5:0] : field_num_1
    ; // @[Serializerhw.scala 115:45 Serializerhw.scala 115:45 Serializerhw.scala 70:28]
  wire [5:0] _GEN_2028 = 4'h2 == stack_num ? class_meta_rsp_fifo_io_out_bits_class_meta_max_field_num[5:0] : field_num_2
    ; // @[Serializerhw.scala 115:45 Serializerhw.scala 115:45 Serializerhw.scala 70:28]
  wire [5:0] _GEN_2029 = 4'h3 == stack_num ? class_meta_rsp_fifo_io_out_bits_class_meta_max_field_num[5:0] : field_num_3
    ; // @[Serializerhw.scala 115:45 Serializerhw.scala 115:45 Serializerhw.scala 70:28]
  wire [5:0] _GEN_2030 = 4'h4 == stack_num ? class_meta_rsp_fifo_io_out_bits_class_meta_max_field_num[5:0] : field_num_4
    ; // @[Serializerhw.scala 115:45 Serializerhw.scala 115:45 Serializerhw.scala 70:28]
  wire [5:0] _GEN_2031 = 4'h5 == stack_num ? class_meta_rsp_fifo_io_out_bits_class_meta_max_field_num[5:0] : field_num_5
    ; // @[Serializerhw.scala 115:45 Serializerhw.scala 115:45 Serializerhw.scala 70:28]
  wire [5:0] _GEN_2032 = 4'h6 == stack_num ? class_meta_rsp_fifo_io_out_bits_class_meta_max_field_num[5:0] : field_num_6
    ; // @[Serializerhw.scala 115:45 Serializerhw.scala 115:45 Serializerhw.scala 70:28]
  wire [5:0] _GEN_2033 = 4'h7 == stack_num ? class_meta_rsp_fifo_io_out_bits_class_meta_max_field_num[5:0] : field_num_7
    ; // @[Serializerhw.scala 115:45 Serializerhw.scala 115:45 Serializerhw.scala 70:28]
  wire [5:0] _GEN_2034 = 4'h8 == stack_num ? class_meta_rsp_fifo_io_out_bits_class_meta_max_field_num[5:0] : field_num_8
    ; // @[Serializerhw.scala 115:45 Serializerhw.scala 115:45 Serializerhw.scala 70:28]
  wire [5:0] _GEN_2035 = 4'h9 == stack_num ? class_meta_rsp_fifo_io_out_bits_class_meta_max_field_num[5:0] : field_num_9
    ; // @[Serializerhw.scala 115:45 Serializerhw.scala 115:45 Serializerhw.scala 70:28]
  wire [5:0] _GEN_2036 = 4'ha == stack_num ? class_meta_rsp_fifo_io_out_bits_class_meta_max_field_num[5:0] :
    field_num_10; // @[Serializerhw.scala 115:45 Serializerhw.scala 115:45 Serializerhw.scala 70:28]
  wire [5:0] _GEN_2037 = 4'hb == stack_num ? class_meta_rsp_fifo_io_out_bits_class_meta_max_field_num[5:0] :
    field_num_11; // @[Serializerhw.scala 115:45 Serializerhw.scala 115:45 Serializerhw.scala 70:28]
  wire [5:0] _GEN_2038 = 4'hc == stack_num ? class_meta_rsp_fifo_io_out_bits_class_meta_max_field_num[5:0] :
    field_num_12; // @[Serializerhw.scala 115:45 Serializerhw.scala 115:45 Serializerhw.scala 70:28]
  wire [5:0] _GEN_2039 = 4'hd == stack_num ? class_meta_rsp_fifo_io_out_bits_class_meta_max_field_num[5:0] :
    field_num_13; // @[Serializerhw.scala 115:45 Serializerhw.scala 115:45 Serializerhw.scala 70:28]
  wire [5:0] _GEN_2040 = 4'he == stack_num ? class_meta_rsp_fifo_io_out_bits_class_meta_max_field_num[5:0] :
    field_num_14; // @[Serializerhw.scala 115:45 Serializerhw.scala 115:45 Serializerhw.scala 70:28]
  wire [5:0] _GEN_2041 = 4'hf == stack_num ? class_meta_rsp_fifo_io_out_bits_class_meta_max_field_num[5:0] :
    field_num_15; // @[Serializerhw.scala 115:45 Serializerhw.scala 115:45 Serializerhw.scala 70:28]
  wire [63:0] _host_base_addr_T_1 = host_base_addr + 64'h400; // @[Serializerhw.scala 117:63]
  wire [7:0] _GEN_4068 = _T_7 ? class_meta_rsp_fifo_io_out_bits_class_meta_max_field_num : {{2'd0}, current_field_num}; // @[Serializerhw.scala 113:52 Serializerhw.scala 116:45 Serializerhw.scala 73:36]
  wire [63:0] _GEN_4071 = _T_7 ? host_base_addr : 64'h0; // @[Serializerhw.scala 113:52 Serializerhw.scala 119:45 Util.scala 13:25]
  wire [31:0] _GEN_4072 = _T_7 ? 32'h40 : 32'h0; // @[Serializerhw.scala 113:52 Serializerhw.scala 120:45 Util.scala 13:25]
  wire  _T_8 = 5'h7 == state; // @[Conditional.scala 37:30]
  wire [4:0] _GEN_4074 = _T_1 ? 5'h13 : state; // @[Serializerhw.scala 125:41 Serializerhw.scala 126:45 Serializerhw.scala 86:46]
  wire  _T_10 = 5'h13 == state; // @[Conditional.scala 37:30]
  wire [4:0] _GEN_4075 = stack_num == 4'h0 ? 5'h10 : 5'he; // @[Serializerhw.scala 131:40 Serializerhw.scala 132:45 Serializerhw.scala 134:45]
  wire  _GEN_10643 = 4'h0 == stack_num; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire  _GEN_10644 = 6'h1 == current_field_num; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4077 = 4'h0 == stack_num & 6'h1 == current_field_num ? field_stack_0_field_type_1_field_type :
    field_stack_0_field_type_0_field_type; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire  _GEN_10646 = 6'h2 == current_field_num; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4078 = 4'h0 == stack_num & 6'h2 == current_field_num ? field_stack_0_field_type_2_field_type :
    _GEN_4077; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire  _GEN_10648 = 6'h3 == current_field_num; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4079 = 4'h0 == stack_num & 6'h3 == current_field_num ? field_stack_0_field_type_3_field_type :
    _GEN_4078; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire  _GEN_10650 = 6'h4 == current_field_num; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4080 = 4'h0 == stack_num & 6'h4 == current_field_num ? field_stack_0_field_type_4_field_type :
    _GEN_4079; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire  _GEN_10652 = 6'h5 == current_field_num; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4081 = 4'h0 == stack_num & 6'h5 == current_field_num ? field_stack_0_field_type_5_field_type :
    _GEN_4080; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire  _GEN_10654 = 6'h6 == current_field_num; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4082 = 4'h0 == stack_num & 6'h6 == current_field_num ? field_stack_0_field_type_6_field_type :
    _GEN_4081; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire  _GEN_10656 = 6'h7 == current_field_num; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4083 = 4'h0 == stack_num & 6'h7 == current_field_num ? field_stack_0_field_type_7_field_type :
    _GEN_4082; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire  _GEN_10658 = 6'h8 == current_field_num; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4084 = 4'h0 == stack_num & 6'h8 == current_field_num ? field_stack_0_field_type_8_field_type :
    _GEN_4083; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire  _GEN_10660 = 6'h9 == current_field_num; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4085 = 4'h0 == stack_num & 6'h9 == current_field_num ? field_stack_0_field_type_9_field_type :
    _GEN_4084; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire  _GEN_10662 = 6'ha == current_field_num; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4086 = 4'h0 == stack_num & 6'ha == current_field_num ? field_stack_0_field_type_10_field_type :
    _GEN_4085; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire  _GEN_10664 = 6'hb == current_field_num; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4087 = 4'h0 == stack_num & 6'hb == current_field_num ? field_stack_0_field_type_11_field_type :
    _GEN_4086; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire  _GEN_10666 = 6'hc == current_field_num; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4088 = 4'h0 == stack_num & 6'hc == current_field_num ? field_stack_0_field_type_12_field_type :
    _GEN_4087; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire  _GEN_10668 = 6'hd == current_field_num; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4089 = 4'h0 == stack_num & 6'hd == current_field_num ? field_stack_0_field_type_13_field_type :
    _GEN_4088; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire  _GEN_10670 = 6'he == current_field_num; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4090 = 4'h0 == stack_num & 6'he == current_field_num ? field_stack_0_field_type_14_field_type :
    _GEN_4089; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire  _GEN_10672 = 6'hf == current_field_num; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4091 = 4'h0 == stack_num & 6'hf == current_field_num ? field_stack_0_field_type_15_field_type :
    _GEN_4090; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire  _GEN_10674 = 6'h10 == current_field_num; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4092 = 4'h0 == stack_num & 6'h10 == current_field_num ? field_stack_0_field_type_16_field_type :
    _GEN_4091; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire  _GEN_10676 = 6'h11 == current_field_num; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4093 = 4'h0 == stack_num & 6'h11 == current_field_num ? field_stack_0_field_type_17_field_type :
    _GEN_4092; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire  _GEN_10678 = 6'h12 == current_field_num; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4094 = 4'h0 == stack_num & 6'h12 == current_field_num ? field_stack_0_field_type_18_field_type :
    _GEN_4093; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire  _GEN_10680 = 6'h13 == current_field_num; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4095 = 4'h0 == stack_num & 6'h13 == current_field_num ? field_stack_0_field_type_19_field_type :
    _GEN_4094; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire  _GEN_10682 = 6'h14 == current_field_num; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4096 = 4'h0 == stack_num & 6'h14 == current_field_num ? field_stack_0_field_type_20_field_type :
    _GEN_4095; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire  _GEN_10684 = 6'h15 == current_field_num; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4097 = 4'h0 == stack_num & 6'h15 == current_field_num ? field_stack_0_field_type_21_field_type :
    _GEN_4096; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire  _GEN_10686 = 6'h16 == current_field_num; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4098 = 4'h0 == stack_num & 6'h16 == current_field_num ? field_stack_0_field_type_22_field_type :
    _GEN_4097; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire  _GEN_10688 = 6'h17 == current_field_num; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4099 = 4'h0 == stack_num & 6'h17 == current_field_num ? field_stack_0_field_type_23_field_type :
    _GEN_4098; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire  _GEN_10690 = 6'h18 == current_field_num; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4100 = 4'h0 == stack_num & 6'h18 == current_field_num ? field_stack_0_field_type_24_field_type :
    _GEN_4099; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire  _GEN_10692 = 6'h19 == current_field_num; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4101 = 4'h0 == stack_num & 6'h19 == current_field_num ? field_stack_0_field_type_25_field_type :
    _GEN_4100; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire  _GEN_10694 = 6'h1a == current_field_num; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4102 = 4'h0 == stack_num & 6'h1a == current_field_num ? field_stack_0_field_type_26_field_type :
    _GEN_4101; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire  _GEN_10696 = 6'h1b == current_field_num; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4103 = 4'h0 == stack_num & 6'h1b == current_field_num ? field_stack_0_field_type_27_field_type :
    _GEN_4102; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire  _GEN_10698 = 6'h1c == current_field_num; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4104 = 4'h0 == stack_num & 6'h1c == current_field_num ? field_stack_0_field_type_28_field_type :
    _GEN_4103; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire  _GEN_10700 = 6'h1d == current_field_num; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4105 = 4'h0 == stack_num & 6'h1d == current_field_num ? field_stack_0_field_type_29_field_type :
    _GEN_4104; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire  _GEN_10702 = 6'h1e == current_field_num; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4106 = 4'h0 == stack_num & 6'h1e == current_field_num ? field_stack_0_field_type_30_field_type :
    _GEN_4105; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire  _GEN_10704 = 6'h1f == current_field_num; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4107 = 4'h0 == stack_num & 6'h1f == current_field_num ? field_stack_0_field_type_31_field_type :
    _GEN_4106; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire  _GEN_10706 = 6'h20 == current_field_num; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4108 = 4'h0 == stack_num & 6'h20 == current_field_num ? field_stack_0_field_type_32_field_type :
    _GEN_4107; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire  _GEN_10707 = 4'h1 == stack_num; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire  _GEN_10708 = 6'h0 == current_field_num; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4109 = 4'h1 == stack_num & 6'h0 == current_field_num ? field_stack_1_field_type_0_field_type :
    _GEN_4108; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4110 = 4'h1 == stack_num & 6'h1 == current_field_num ? field_stack_1_field_type_1_field_type :
    _GEN_4109; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4111 = 4'h1 == stack_num & 6'h2 == current_field_num ? field_stack_1_field_type_2_field_type :
    _GEN_4110; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4112 = 4'h1 == stack_num & 6'h3 == current_field_num ? field_stack_1_field_type_3_field_type :
    _GEN_4111; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4113 = 4'h1 == stack_num & 6'h4 == current_field_num ? field_stack_1_field_type_4_field_type :
    _GEN_4112; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4114 = 4'h1 == stack_num & 6'h5 == current_field_num ? field_stack_1_field_type_5_field_type :
    _GEN_4113; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4115 = 4'h1 == stack_num & 6'h6 == current_field_num ? field_stack_1_field_type_6_field_type :
    _GEN_4114; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4116 = 4'h1 == stack_num & 6'h7 == current_field_num ? field_stack_1_field_type_7_field_type :
    _GEN_4115; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4117 = 4'h1 == stack_num & 6'h8 == current_field_num ? field_stack_1_field_type_8_field_type :
    _GEN_4116; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4118 = 4'h1 == stack_num & 6'h9 == current_field_num ? field_stack_1_field_type_9_field_type :
    _GEN_4117; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4119 = 4'h1 == stack_num & 6'ha == current_field_num ? field_stack_1_field_type_10_field_type :
    _GEN_4118; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4120 = 4'h1 == stack_num & 6'hb == current_field_num ? field_stack_1_field_type_11_field_type :
    _GEN_4119; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4121 = 4'h1 == stack_num & 6'hc == current_field_num ? field_stack_1_field_type_12_field_type :
    _GEN_4120; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4122 = 4'h1 == stack_num & 6'hd == current_field_num ? field_stack_1_field_type_13_field_type :
    _GEN_4121; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4123 = 4'h1 == stack_num & 6'he == current_field_num ? field_stack_1_field_type_14_field_type :
    _GEN_4122; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4124 = 4'h1 == stack_num & 6'hf == current_field_num ? field_stack_1_field_type_15_field_type :
    _GEN_4123; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4125 = 4'h1 == stack_num & 6'h10 == current_field_num ? field_stack_1_field_type_16_field_type :
    _GEN_4124; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4126 = 4'h1 == stack_num & 6'h11 == current_field_num ? field_stack_1_field_type_17_field_type :
    _GEN_4125; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4127 = 4'h1 == stack_num & 6'h12 == current_field_num ? field_stack_1_field_type_18_field_type :
    _GEN_4126; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4128 = 4'h1 == stack_num & 6'h13 == current_field_num ? field_stack_1_field_type_19_field_type :
    _GEN_4127; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4129 = 4'h1 == stack_num & 6'h14 == current_field_num ? field_stack_1_field_type_20_field_type :
    _GEN_4128; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4130 = 4'h1 == stack_num & 6'h15 == current_field_num ? field_stack_1_field_type_21_field_type :
    _GEN_4129; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4131 = 4'h1 == stack_num & 6'h16 == current_field_num ? field_stack_1_field_type_22_field_type :
    _GEN_4130; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4132 = 4'h1 == stack_num & 6'h17 == current_field_num ? field_stack_1_field_type_23_field_type :
    _GEN_4131; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4133 = 4'h1 == stack_num & 6'h18 == current_field_num ? field_stack_1_field_type_24_field_type :
    _GEN_4132; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4134 = 4'h1 == stack_num & 6'h19 == current_field_num ? field_stack_1_field_type_25_field_type :
    _GEN_4133; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4135 = 4'h1 == stack_num & 6'h1a == current_field_num ? field_stack_1_field_type_26_field_type :
    _GEN_4134; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4136 = 4'h1 == stack_num & 6'h1b == current_field_num ? field_stack_1_field_type_27_field_type :
    _GEN_4135; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4137 = 4'h1 == stack_num & 6'h1c == current_field_num ? field_stack_1_field_type_28_field_type :
    _GEN_4136; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4138 = 4'h1 == stack_num & 6'h1d == current_field_num ? field_stack_1_field_type_29_field_type :
    _GEN_4137; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4139 = 4'h1 == stack_num & 6'h1e == current_field_num ? field_stack_1_field_type_30_field_type :
    _GEN_4138; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4140 = 4'h1 == stack_num & 6'h1f == current_field_num ? field_stack_1_field_type_31_field_type :
    _GEN_4139; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4141 = 4'h1 == stack_num & 6'h20 == current_field_num ? field_stack_1_field_type_32_field_type :
    _GEN_4140; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire  _GEN_10773 = 4'h2 == stack_num; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4142 = 4'h2 == stack_num & 6'h0 == current_field_num ? field_stack_2_field_type_0_field_type :
    _GEN_4141; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4143 = 4'h2 == stack_num & 6'h1 == current_field_num ? field_stack_2_field_type_1_field_type :
    _GEN_4142; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4144 = 4'h2 == stack_num & 6'h2 == current_field_num ? field_stack_2_field_type_2_field_type :
    _GEN_4143; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4145 = 4'h2 == stack_num & 6'h3 == current_field_num ? field_stack_2_field_type_3_field_type :
    _GEN_4144; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4146 = 4'h2 == stack_num & 6'h4 == current_field_num ? field_stack_2_field_type_4_field_type :
    _GEN_4145; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4147 = 4'h2 == stack_num & 6'h5 == current_field_num ? field_stack_2_field_type_5_field_type :
    _GEN_4146; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4148 = 4'h2 == stack_num & 6'h6 == current_field_num ? field_stack_2_field_type_6_field_type :
    _GEN_4147; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4149 = 4'h2 == stack_num & 6'h7 == current_field_num ? field_stack_2_field_type_7_field_type :
    _GEN_4148; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4150 = 4'h2 == stack_num & 6'h8 == current_field_num ? field_stack_2_field_type_8_field_type :
    _GEN_4149; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4151 = 4'h2 == stack_num & 6'h9 == current_field_num ? field_stack_2_field_type_9_field_type :
    _GEN_4150; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4152 = 4'h2 == stack_num & 6'ha == current_field_num ? field_stack_2_field_type_10_field_type :
    _GEN_4151; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4153 = 4'h2 == stack_num & 6'hb == current_field_num ? field_stack_2_field_type_11_field_type :
    _GEN_4152; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4154 = 4'h2 == stack_num & 6'hc == current_field_num ? field_stack_2_field_type_12_field_type :
    _GEN_4153; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4155 = 4'h2 == stack_num & 6'hd == current_field_num ? field_stack_2_field_type_13_field_type :
    _GEN_4154; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4156 = 4'h2 == stack_num & 6'he == current_field_num ? field_stack_2_field_type_14_field_type :
    _GEN_4155; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4157 = 4'h2 == stack_num & 6'hf == current_field_num ? field_stack_2_field_type_15_field_type :
    _GEN_4156; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4158 = 4'h2 == stack_num & 6'h10 == current_field_num ? field_stack_2_field_type_16_field_type :
    _GEN_4157; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4159 = 4'h2 == stack_num & 6'h11 == current_field_num ? field_stack_2_field_type_17_field_type :
    _GEN_4158; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4160 = 4'h2 == stack_num & 6'h12 == current_field_num ? field_stack_2_field_type_18_field_type :
    _GEN_4159; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4161 = 4'h2 == stack_num & 6'h13 == current_field_num ? field_stack_2_field_type_19_field_type :
    _GEN_4160; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4162 = 4'h2 == stack_num & 6'h14 == current_field_num ? field_stack_2_field_type_20_field_type :
    _GEN_4161; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4163 = 4'h2 == stack_num & 6'h15 == current_field_num ? field_stack_2_field_type_21_field_type :
    _GEN_4162; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4164 = 4'h2 == stack_num & 6'h16 == current_field_num ? field_stack_2_field_type_22_field_type :
    _GEN_4163; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4165 = 4'h2 == stack_num & 6'h17 == current_field_num ? field_stack_2_field_type_23_field_type :
    _GEN_4164; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4166 = 4'h2 == stack_num & 6'h18 == current_field_num ? field_stack_2_field_type_24_field_type :
    _GEN_4165; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4167 = 4'h2 == stack_num & 6'h19 == current_field_num ? field_stack_2_field_type_25_field_type :
    _GEN_4166; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4168 = 4'h2 == stack_num & 6'h1a == current_field_num ? field_stack_2_field_type_26_field_type :
    _GEN_4167; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4169 = 4'h2 == stack_num & 6'h1b == current_field_num ? field_stack_2_field_type_27_field_type :
    _GEN_4168; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4170 = 4'h2 == stack_num & 6'h1c == current_field_num ? field_stack_2_field_type_28_field_type :
    _GEN_4169; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4171 = 4'h2 == stack_num & 6'h1d == current_field_num ? field_stack_2_field_type_29_field_type :
    _GEN_4170; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4172 = 4'h2 == stack_num & 6'h1e == current_field_num ? field_stack_2_field_type_30_field_type :
    _GEN_4171; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4173 = 4'h2 == stack_num & 6'h1f == current_field_num ? field_stack_2_field_type_31_field_type :
    _GEN_4172; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4174 = 4'h2 == stack_num & 6'h20 == current_field_num ? field_stack_2_field_type_32_field_type :
    _GEN_4173; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire  _GEN_10839 = 4'h3 == stack_num; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4175 = 4'h3 == stack_num & 6'h0 == current_field_num ? field_stack_3_field_type_0_field_type :
    _GEN_4174; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4176 = 4'h3 == stack_num & 6'h1 == current_field_num ? field_stack_3_field_type_1_field_type :
    _GEN_4175; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4177 = 4'h3 == stack_num & 6'h2 == current_field_num ? field_stack_3_field_type_2_field_type :
    _GEN_4176; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4178 = 4'h3 == stack_num & 6'h3 == current_field_num ? field_stack_3_field_type_3_field_type :
    _GEN_4177; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4179 = 4'h3 == stack_num & 6'h4 == current_field_num ? field_stack_3_field_type_4_field_type :
    _GEN_4178; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4180 = 4'h3 == stack_num & 6'h5 == current_field_num ? field_stack_3_field_type_5_field_type :
    _GEN_4179; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4181 = 4'h3 == stack_num & 6'h6 == current_field_num ? field_stack_3_field_type_6_field_type :
    _GEN_4180; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4182 = 4'h3 == stack_num & 6'h7 == current_field_num ? field_stack_3_field_type_7_field_type :
    _GEN_4181; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4183 = 4'h3 == stack_num & 6'h8 == current_field_num ? field_stack_3_field_type_8_field_type :
    _GEN_4182; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4184 = 4'h3 == stack_num & 6'h9 == current_field_num ? field_stack_3_field_type_9_field_type :
    _GEN_4183; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4185 = 4'h3 == stack_num & 6'ha == current_field_num ? field_stack_3_field_type_10_field_type :
    _GEN_4184; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4186 = 4'h3 == stack_num & 6'hb == current_field_num ? field_stack_3_field_type_11_field_type :
    _GEN_4185; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4187 = 4'h3 == stack_num & 6'hc == current_field_num ? field_stack_3_field_type_12_field_type :
    _GEN_4186; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4188 = 4'h3 == stack_num & 6'hd == current_field_num ? field_stack_3_field_type_13_field_type :
    _GEN_4187; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4189 = 4'h3 == stack_num & 6'he == current_field_num ? field_stack_3_field_type_14_field_type :
    _GEN_4188; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4190 = 4'h3 == stack_num & 6'hf == current_field_num ? field_stack_3_field_type_15_field_type :
    _GEN_4189; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4191 = 4'h3 == stack_num & 6'h10 == current_field_num ? field_stack_3_field_type_16_field_type :
    _GEN_4190; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4192 = 4'h3 == stack_num & 6'h11 == current_field_num ? field_stack_3_field_type_17_field_type :
    _GEN_4191; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4193 = 4'h3 == stack_num & 6'h12 == current_field_num ? field_stack_3_field_type_18_field_type :
    _GEN_4192; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4194 = 4'h3 == stack_num & 6'h13 == current_field_num ? field_stack_3_field_type_19_field_type :
    _GEN_4193; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4195 = 4'h3 == stack_num & 6'h14 == current_field_num ? field_stack_3_field_type_20_field_type :
    _GEN_4194; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4196 = 4'h3 == stack_num & 6'h15 == current_field_num ? field_stack_3_field_type_21_field_type :
    _GEN_4195; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4197 = 4'h3 == stack_num & 6'h16 == current_field_num ? field_stack_3_field_type_22_field_type :
    _GEN_4196; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4198 = 4'h3 == stack_num & 6'h17 == current_field_num ? field_stack_3_field_type_23_field_type :
    _GEN_4197; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4199 = 4'h3 == stack_num & 6'h18 == current_field_num ? field_stack_3_field_type_24_field_type :
    _GEN_4198; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4200 = 4'h3 == stack_num & 6'h19 == current_field_num ? field_stack_3_field_type_25_field_type :
    _GEN_4199; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4201 = 4'h3 == stack_num & 6'h1a == current_field_num ? field_stack_3_field_type_26_field_type :
    _GEN_4200; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4202 = 4'h3 == stack_num & 6'h1b == current_field_num ? field_stack_3_field_type_27_field_type :
    _GEN_4201; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4203 = 4'h3 == stack_num & 6'h1c == current_field_num ? field_stack_3_field_type_28_field_type :
    _GEN_4202; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4204 = 4'h3 == stack_num & 6'h1d == current_field_num ? field_stack_3_field_type_29_field_type :
    _GEN_4203; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4205 = 4'h3 == stack_num & 6'h1e == current_field_num ? field_stack_3_field_type_30_field_type :
    _GEN_4204; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4206 = 4'h3 == stack_num & 6'h1f == current_field_num ? field_stack_3_field_type_31_field_type :
    _GEN_4205; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4207 = 4'h3 == stack_num & 6'h20 == current_field_num ? field_stack_3_field_type_32_field_type :
    _GEN_4206; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire  _GEN_10905 = 4'h4 == stack_num; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4208 = 4'h4 == stack_num & 6'h0 == current_field_num ? field_stack_4_field_type_0_field_type :
    _GEN_4207; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4209 = 4'h4 == stack_num & 6'h1 == current_field_num ? field_stack_4_field_type_1_field_type :
    _GEN_4208; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4210 = 4'h4 == stack_num & 6'h2 == current_field_num ? field_stack_4_field_type_2_field_type :
    _GEN_4209; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4211 = 4'h4 == stack_num & 6'h3 == current_field_num ? field_stack_4_field_type_3_field_type :
    _GEN_4210; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4212 = 4'h4 == stack_num & 6'h4 == current_field_num ? field_stack_4_field_type_4_field_type :
    _GEN_4211; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4213 = 4'h4 == stack_num & 6'h5 == current_field_num ? field_stack_4_field_type_5_field_type :
    _GEN_4212; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4214 = 4'h4 == stack_num & 6'h6 == current_field_num ? field_stack_4_field_type_6_field_type :
    _GEN_4213; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4215 = 4'h4 == stack_num & 6'h7 == current_field_num ? field_stack_4_field_type_7_field_type :
    _GEN_4214; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4216 = 4'h4 == stack_num & 6'h8 == current_field_num ? field_stack_4_field_type_8_field_type :
    _GEN_4215; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4217 = 4'h4 == stack_num & 6'h9 == current_field_num ? field_stack_4_field_type_9_field_type :
    _GEN_4216; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4218 = 4'h4 == stack_num & 6'ha == current_field_num ? field_stack_4_field_type_10_field_type :
    _GEN_4217; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4219 = 4'h4 == stack_num & 6'hb == current_field_num ? field_stack_4_field_type_11_field_type :
    _GEN_4218; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4220 = 4'h4 == stack_num & 6'hc == current_field_num ? field_stack_4_field_type_12_field_type :
    _GEN_4219; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4221 = 4'h4 == stack_num & 6'hd == current_field_num ? field_stack_4_field_type_13_field_type :
    _GEN_4220; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4222 = 4'h4 == stack_num & 6'he == current_field_num ? field_stack_4_field_type_14_field_type :
    _GEN_4221; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4223 = 4'h4 == stack_num & 6'hf == current_field_num ? field_stack_4_field_type_15_field_type :
    _GEN_4222; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4224 = 4'h4 == stack_num & 6'h10 == current_field_num ? field_stack_4_field_type_16_field_type :
    _GEN_4223; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4225 = 4'h4 == stack_num & 6'h11 == current_field_num ? field_stack_4_field_type_17_field_type :
    _GEN_4224; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4226 = 4'h4 == stack_num & 6'h12 == current_field_num ? field_stack_4_field_type_18_field_type :
    _GEN_4225; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4227 = 4'h4 == stack_num & 6'h13 == current_field_num ? field_stack_4_field_type_19_field_type :
    _GEN_4226; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4228 = 4'h4 == stack_num & 6'h14 == current_field_num ? field_stack_4_field_type_20_field_type :
    _GEN_4227; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4229 = 4'h4 == stack_num & 6'h15 == current_field_num ? field_stack_4_field_type_21_field_type :
    _GEN_4228; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4230 = 4'h4 == stack_num & 6'h16 == current_field_num ? field_stack_4_field_type_22_field_type :
    _GEN_4229; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4231 = 4'h4 == stack_num & 6'h17 == current_field_num ? field_stack_4_field_type_23_field_type :
    _GEN_4230; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4232 = 4'h4 == stack_num & 6'h18 == current_field_num ? field_stack_4_field_type_24_field_type :
    _GEN_4231; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4233 = 4'h4 == stack_num & 6'h19 == current_field_num ? field_stack_4_field_type_25_field_type :
    _GEN_4232; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4234 = 4'h4 == stack_num & 6'h1a == current_field_num ? field_stack_4_field_type_26_field_type :
    _GEN_4233; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4235 = 4'h4 == stack_num & 6'h1b == current_field_num ? field_stack_4_field_type_27_field_type :
    _GEN_4234; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4236 = 4'h4 == stack_num & 6'h1c == current_field_num ? field_stack_4_field_type_28_field_type :
    _GEN_4235; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4237 = 4'h4 == stack_num & 6'h1d == current_field_num ? field_stack_4_field_type_29_field_type :
    _GEN_4236; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4238 = 4'h4 == stack_num & 6'h1e == current_field_num ? field_stack_4_field_type_30_field_type :
    _GEN_4237; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4239 = 4'h4 == stack_num & 6'h1f == current_field_num ? field_stack_4_field_type_31_field_type :
    _GEN_4238; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4240 = 4'h4 == stack_num & 6'h20 == current_field_num ? field_stack_4_field_type_32_field_type :
    _GEN_4239; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire  _GEN_10971 = 4'h5 == stack_num; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4241 = 4'h5 == stack_num & 6'h0 == current_field_num ? field_stack_5_field_type_0_field_type :
    _GEN_4240; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4242 = 4'h5 == stack_num & 6'h1 == current_field_num ? field_stack_5_field_type_1_field_type :
    _GEN_4241; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4243 = 4'h5 == stack_num & 6'h2 == current_field_num ? field_stack_5_field_type_2_field_type :
    _GEN_4242; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4244 = 4'h5 == stack_num & 6'h3 == current_field_num ? field_stack_5_field_type_3_field_type :
    _GEN_4243; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4245 = 4'h5 == stack_num & 6'h4 == current_field_num ? field_stack_5_field_type_4_field_type :
    _GEN_4244; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4246 = 4'h5 == stack_num & 6'h5 == current_field_num ? field_stack_5_field_type_5_field_type :
    _GEN_4245; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4247 = 4'h5 == stack_num & 6'h6 == current_field_num ? field_stack_5_field_type_6_field_type :
    _GEN_4246; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4248 = 4'h5 == stack_num & 6'h7 == current_field_num ? field_stack_5_field_type_7_field_type :
    _GEN_4247; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4249 = 4'h5 == stack_num & 6'h8 == current_field_num ? field_stack_5_field_type_8_field_type :
    _GEN_4248; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4250 = 4'h5 == stack_num & 6'h9 == current_field_num ? field_stack_5_field_type_9_field_type :
    _GEN_4249; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4251 = 4'h5 == stack_num & 6'ha == current_field_num ? field_stack_5_field_type_10_field_type :
    _GEN_4250; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4252 = 4'h5 == stack_num & 6'hb == current_field_num ? field_stack_5_field_type_11_field_type :
    _GEN_4251; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4253 = 4'h5 == stack_num & 6'hc == current_field_num ? field_stack_5_field_type_12_field_type :
    _GEN_4252; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4254 = 4'h5 == stack_num & 6'hd == current_field_num ? field_stack_5_field_type_13_field_type :
    _GEN_4253; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4255 = 4'h5 == stack_num & 6'he == current_field_num ? field_stack_5_field_type_14_field_type :
    _GEN_4254; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4256 = 4'h5 == stack_num & 6'hf == current_field_num ? field_stack_5_field_type_15_field_type :
    _GEN_4255; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4257 = 4'h5 == stack_num & 6'h10 == current_field_num ? field_stack_5_field_type_16_field_type :
    _GEN_4256; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4258 = 4'h5 == stack_num & 6'h11 == current_field_num ? field_stack_5_field_type_17_field_type :
    _GEN_4257; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4259 = 4'h5 == stack_num & 6'h12 == current_field_num ? field_stack_5_field_type_18_field_type :
    _GEN_4258; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4260 = 4'h5 == stack_num & 6'h13 == current_field_num ? field_stack_5_field_type_19_field_type :
    _GEN_4259; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4261 = 4'h5 == stack_num & 6'h14 == current_field_num ? field_stack_5_field_type_20_field_type :
    _GEN_4260; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4262 = 4'h5 == stack_num & 6'h15 == current_field_num ? field_stack_5_field_type_21_field_type :
    _GEN_4261; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4263 = 4'h5 == stack_num & 6'h16 == current_field_num ? field_stack_5_field_type_22_field_type :
    _GEN_4262; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4264 = 4'h5 == stack_num & 6'h17 == current_field_num ? field_stack_5_field_type_23_field_type :
    _GEN_4263; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4265 = 4'h5 == stack_num & 6'h18 == current_field_num ? field_stack_5_field_type_24_field_type :
    _GEN_4264; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4266 = 4'h5 == stack_num & 6'h19 == current_field_num ? field_stack_5_field_type_25_field_type :
    _GEN_4265; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4267 = 4'h5 == stack_num & 6'h1a == current_field_num ? field_stack_5_field_type_26_field_type :
    _GEN_4266; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4268 = 4'h5 == stack_num & 6'h1b == current_field_num ? field_stack_5_field_type_27_field_type :
    _GEN_4267; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4269 = 4'h5 == stack_num & 6'h1c == current_field_num ? field_stack_5_field_type_28_field_type :
    _GEN_4268; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4270 = 4'h5 == stack_num & 6'h1d == current_field_num ? field_stack_5_field_type_29_field_type :
    _GEN_4269; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4271 = 4'h5 == stack_num & 6'h1e == current_field_num ? field_stack_5_field_type_30_field_type :
    _GEN_4270; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4272 = 4'h5 == stack_num & 6'h1f == current_field_num ? field_stack_5_field_type_31_field_type :
    _GEN_4271; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4273 = 4'h5 == stack_num & 6'h20 == current_field_num ? field_stack_5_field_type_32_field_type :
    _GEN_4272; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire  _GEN_11037 = 4'h6 == stack_num; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4274 = 4'h6 == stack_num & 6'h0 == current_field_num ? field_stack_6_field_type_0_field_type :
    _GEN_4273; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4275 = 4'h6 == stack_num & 6'h1 == current_field_num ? field_stack_6_field_type_1_field_type :
    _GEN_4274; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4276 = 4'h6 == stack_num & 6'h2 == current_field_num ? field_stack_6_field_type_2_field_type :
    _GEN_4275; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4277 = 4'h6 == stack_num & 6'h3 == current_field_num ? field_stack_6_field_type_3_field_type :
    _GEN_4276; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4278 = 4'h6 == stack_num & 6'h4 == current_field_num ? field_stack_6_field_type_4_field_type :
    _GEN_4277; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4279 = 4'h6 == stack_num & 6'h5 == current_field_num ? field_stack_6_field_type_5_field_type :
    _GEN_4278; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4280 = 4'h6 == stack_num & 6'h6 == current_field_num ? field_stack_6_field_type_6_field_type :
    _GEN_4279; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4281 = 4'h6 == stack_num & 6'h7 == current_field_num ? field_stack_6_field_type_7_field_type :
    _GEN_4280; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4282 = 4'h6 == stack_num & 6'h8 == current_field_num ? field_stack_6_field_type_8_field_type :
    _GEN_4281; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4283 = 4'h6 == stack_num & 6'h9 == current_field_num ? field_stack_6_field_type_9_field_type :
    _GEN_4282; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4284 = 4'h6 == stack_num & 6'ha == current_field_num ? field_stack_6_field_type_10_field_type :
    _GEN_4283; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4285 = 4'h6 == stack_num & 6'hb == current_field_num ? field_stack_6_field_type_11_field_type :
    _GEN_4284; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4286 = 4'h6 == stack_num & 6'hc == current_field_num ? field_stack_6_field_type_12_field_type :
    _GEN_4285; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4287 = 4'h6 == stack_num & 6'hd == current_field_num ? field_stack_6_field_type_13_field_type :
    _GEN_4286; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4288 = 4'h6 == stack_num & 6'he == current_field_num ? field_stack_6_field_type_14_field_type :
    _GEN_4287; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4289 = 4'h6 == stack_num & 6'hf == current_field_num ? field_stack_6_field_type_15_field_type :
    _GEN_4288; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4290 = 4'h6 == stack_num & 6'h10 == current_field_num ? field_stack_6_field_type_16_field_type :
    _GEN_4289; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4291 = 4'h6 == stack_num & 6'h11 == current_field_num ? field_stack_6_field_type_17_field_type :
    _GEN_4290; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4292 = 4'h6 == stack_num & 6'h12 == current_field_num ? field_stack_6_field_type_18_field_type :
    _GEN_4291; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4293 = 4'h6 == stack_num & 6'h13 == current_field_num ? field_stack_6_field_type_19_field_type :
    _GEN_4292; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4294 = 4'h6 == stack_num & 6'h14 == current_field_num ? field_stack_6_field_type_20_field_type :
    _GEN_4293; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4295 = 4'h6 == stack_num & 6'h15 == current_field_num ? field_stack_6_field_type_21_field_type :
    _GEN_4294; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4296 = 4'h6 == stack_num & 6'h16 == current_field_num ? field_stack_6_field_type_22_field_type :
    _GEN_4295; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4297 = 4'h6 == stack_num & 6'h17 == current_field_num ? field_stack_6_field_type_23_field_type :
    _GEN_4296; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4298 = 4'h6 == stack_num & 6'h18 == current_field_num ? field_stack_6_field_type_24_field_type :
    _GEN_4297; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4299 = 4'h6 == stack_num & 6'h19 == current_field_num ? field_stack_6_field_type_25_field_type :
    _GEN_4298; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4300 = 4'h6 == stack_num & 6'h1a == current_field_num ? field_stack_6_field_type_26_field_type :
    _GEN_4299; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4301 = 4'h6 == stack_num & 6'h1b == current_field_num ? field_stack_6_field_type_27_field_type :
    _GEN_4300; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4302 = 4'h6 == stack_num & 6'h1c == current_field_num ? field_stack_6_field_type_28_field_type :
    _GEN_4301; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4303 = 4'h6 == stack_num & 6'h1d == current_field_num ? field_stack_6_field_type_29_field_type :
    _GEN_4302; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4304 = 4'h6 == stack_num & 6'h1e == current_field_num ? field_stack_6_field_type_30_field_type :
    _GEN_4303; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4305 = 4'h6 == stack_num & 6'h1f == current_field_num ? field_stack_6_field_type_31_field_type :
    _GEN_4304; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4306 = 4'h6 == stack_num & 6'h20 == current_field_num ? field_stack_6_field_type_32_field_type :
    _GEN_4305; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire  _GEN_11103 = 4'h7 == stack_num; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4307 = 4'h7 == stack_num & 6'h0 == current_field_num ? field_stack_7_field_type_0_field_type :
    _GEN_4306; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4308 = 4'h7 == stack_num & 6'h1 == current_field_num ? field_stack_7_field_type_1_field_type :
    _GEN_4307; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4309 = 4'h7 == stack_num & 6'h2 == current_field_num ? field_stack_7_field_type_2_field_type :
    _GEN_4308; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4310 = 4'h7 == stack_num & 6'h3 == current_field_num ? field_stack_7_field_type_3_field_type :
    _GEN_4309; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4311 = 4'h7 == stack_num & 6'h4 == current_field_num ? field_stack_7_field_type_4_field_type :
    _GEN_4310; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4312 = 4'h7 == stack_num & 6'h5 == current_field_num ? field_stack_7_field_type_5_field_type :
    _GEN_4311; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4313 = 4'h7 == stack_num & 6'h6 == current_field_num ? field_stack_7_field_type_6_field_type :
    _GEN_4312; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4314 = 4'h7 == stack_num & 6'h7 == current_field_num ? field_stack_7_field_type_7_field_type :
    _GEN_4313; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4315 = 4'h7 == stack_num & 6'h8 == current_field_num ? field_stack_7_field_type_8_field_type :
    _GEN_4314; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4316 = 4'h7 == stack_num & 6'h9 == current_field_num ? field_stack_7_field_type_9_field_type :
    _GEN_4315; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4317 = 4'h7 == stack_num & 6'ha == current_field_num ? field_stack_7_field_type_10_field_type :
    _GEN_4316; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4318 = 4'h7 == stack_num & 6'hb == current_field_num ? field_stack_7_field_type_11_field_type :
    _GEN_4317; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4319 = 4'h7 == stack_num & 6'hc == current_field_num ? field_stack_7_field_type_12_field_type :
    _GEN_4318; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4320 = 4'h7 == stack_num & 6'hd == current_field_num ? field_stack_7_field_type_13_field_type :
    _GEN_4319; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4321 = 4'h7 == stack_num & 6'he == current_field_num ? field_stack_7_field_type_14_field_type :
    _GEN_4320; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4322 = 4'h7 == stack_num & 6'hf == current_field_num ? field_stack_7_field_type_15_field_type :
    _GEN_4321; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4323 = 4'h7 == stack_num & 6'h10 == current_field_num ? field_stack_7_field_type_16_field_type :
    _GEN_4322; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4324 = 4'h7 == stack_num & 6'h11 == current_field_num ? field_stack_7_field_type_17_field_type :
    _GEN_4323; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4325 = 4'h7 == stack_num & 6'h12 == current_field_num ? field_stack_7_field_type_18_field_type :
    _GEN_4324; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4326 = 4'h7 == stack_num & 6'h13 == current_field_num ? field_stack_7_field_type_19_field_type :
    _GEN_4325; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4327 = 4'h7 == stack_num & 6'h14 == current_field_num ? field_stack_7_field_type_20_field_type :
    _GEN_4326; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4328 = 4'h7 == stack_num & 6'h15 == current_field_num ? field_stack_7_field_type_21_field_type :
    _GEN_4327; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4329 = 4'h7 == stack_num & 6'h16 == current_field_num ? field_stack_7_field_type_22_field_type :
    _GEN_4328; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4330 = 4'h7 == stack_num & 6'h17 == current_field_num ? field_stack_7_field_type_23_field_type :
    _GEN_4329; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4331 = 4'h7 == stack_num & 6'h18 == current_field_num ? field_stack_7_field_type_24_field_type :
    _GEN_4330; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4332 = 4'h7 == stack_num & 6'h19 == current_field_num ? field_stack_7_field_type_25_field_type :
    _GEN_4331; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4333 = 4'h7 == stack_num & 6'h1a == current_field_num ? field_stack_7_field_type_26_field_type :
    _GEN_4332; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4334 = 4'h7 == stack_num & 6'h1b == current_field_num ? field_stack_7_field_type_27_field_type :
    _GEN_4333; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4335 = 4'h7 == stack_num & 6'h1c == current_field_num ? field_stack_7_field_type_28_field_type :
    _GEN_4334; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4336 = 4'h7 == stack_num & 6'h1d == current_field_num ? field_stack_7_field_type_29_field_type :
    _GEN_4335; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4337 = 4'h7 == stack_num & 6'h1e == current_field_num ? field_stack_7_field_type_30_field_type :
    _GEN_4336; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4338 = 4'h7 == stack_num & 6'h1f == current_field_num ? field_stack_7_field_type_31_field_type :
    _GEN_4337; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4339 = 4'h7 == stack_num & 6'h20 == current_field_num ? field_stack_7_field_type_32_field_type :
    _GEN_4338; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire  _GEN_11169 = 4'h8 == stack_num; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4340 = 4'h8 == stack_num & 6'h0 == current_field_num ? field_stack_8_field_type_0_field_type :
    _GEN_4339; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4341 = 4'h8 == stack_num & 6'h1 == current_field_num ? field_stack_8_field_type_1_field_type :
    _GEN_4340; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4342 = 4'h8 == stack_num & 6'h2 == current_field_num ? field_stack_8_field_type_2_field_type :
    _GEN_4341; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4343 = 4'h8 == stack_num & 6'h3 == current_field_num ? field_stack_8_field_type_3_field_type :
    _GEN_4342; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4344 = 4'h8 == stack_num & 6'h4 == current_field_num ? field_stack_8_field_type_4_field_type :
    _GEN_4343; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4345 = 4'h8 == stack_num & 6'h5 == current_field_num ? field_stack_8_field_type_5_field_type :
    _GEN_4344; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4346 = 4'h8 == stack_num & 6'h6 == current_field_num ? field_stack_8_field_type_6_field_type :
    _GEN_4345; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4347 = 4'h8 == stack_num & 6'h7 == current_field_num ? field_stack_8_field_type_7_field_type :
    _GEN_4346; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4348 = 4'h8 == stack_num & 6'h8 == current_field_num ? field_stack_8_field_type_8_field_type :
    _GEN_4347; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4349 = 4'h8 == stack_num & 6'h9 == current_field_num ? field_stack_8_field_type_9_field_type :
    _GEN_4348; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4350 = 4'h8 == stack_num & 6'ha == current_field_num ? field_stack_8_field_type_10_field_type :
    _GEN_4349; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4351 = 4'h8 == stack_num & 6'hb == current_field_num ? field_stack_8_field_type_11_field_type :
    _GEN_4350; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4352 = 4'h8 == stack_num & 6'hc == current_field_num ? field_stack_8_field_type_12_field_type :
    _GEN_4351; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4353 = 4'h8 == stack_num & 6'hd == current_field_num ? field_stack_8_field_type_13_field_type :
    _GEN_4352; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4354 = 4'h8 == stack_num & 6'he == current_field_num ? field_stack_8_field_type_14_field_type :
    _GEN_4353; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4355 = 4'h8 == stack_num & 6'hf == current_field_num ? field_stack_8_field_type_15_field_type :
    _GEN_4354; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4356 = 4'h8 == stack_num & 6'h10 == current_field_num ? field_stack_8_field_type_16_field_type :
    _GEN_4355; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4357 = 4'h8 == stack_num & 6'h11 == current_field_num ? field_stack_8_field_type_17_field_type :
    _GEN_4356; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4358 = 4'h8 == stack_num & 6'h12 == current_field_num ? field_stack_8_field_type_18_field_type :
    _GEN_4357; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4359 = 4'h8 == stack_num & 6'h13 == current_field_num ? field_stack_8_field_type_19_field_type :
    _GEN_4358; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4360 = 4'h8 == stack_num & 6'h14 == current_field_num ? field_stack_8_field_type_20_field_type :
    _GEN_4359; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4361 = 4'h8 == stack_num & 6'h15 == current_field_num ? field_stack_8_field_type_21_field_type :
    _GEN_4360; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4362 = 4'h8 == stack_num & 6'h16 == current_field_num ? field_stack_8_field_type_22_field_type :
    _GEN_4361; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4363 = 4'h8 == stack_num & 6'h17 == current_field_num ? field_stack_8_field_type_23_field_type :
    _GEN_4362; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4364 = 4'h8 == stack_num & 6'h18 == current_field_num ? field_stack_8_field_type_24_field_type :
    _GEN_4363; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4365 = 4'h8 == stack_num & 6'h19 == current_field_num ? field_stack_8_field_type_25_field_type :
    _GEN_4364; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4366 = 4'h8 == stack_num & 6'h1a == current_field_num ? field_stack_8_field_type_26_field_type :
    _GEN_4365; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4367 = 4'h8 == stack_num & 6'h1b == current_field_num ? field_stack_8_field_type_27_field_type :
    _GEN_4366; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4368 = 4'h8 == stack_num & 6'h1c == current_field_num ? field_stack_8_field_type_28_field_type :
    _GEN_4367; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4369 = 4'h8 == stack_num & 6'h1d == current_field_num ? field_stack_8_field_type_29_field_type :
    _GEN_4368; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4370 = 4'h8 == stack_num & 6'h1e == current_field_num ? field_stack_8_field_type_30_field_type :
    _GEN_4369; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4371 = 4'h8 == stack_num & 6'h1f == current_field_num ? field_stack_8_field_type_31_field_type :
    _GEN_4370; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4372 = 4'h8 == stack_num & 6'h20 == current_field_num ? field_stack_8_field_type_32_field_type :
    _GEN_4371; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire  _GEN_11235 = 4'h9 == stack_num; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4373 = 4'h9 == stack_num & 6'h0 == current_field_num ? field_stack_9_field_type_0_field_type :
    _GEN_4372; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4374 = 4'h9 == stack_num & 6'h1 == current_field_num ? field_stack_9_field_type_1_field_type :
    _GEN_4373; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4375 = 4'h9 == stack_num & 6'h2 == current_field_num ? field_stack_9_field_type_2_field_type :
    _GEN_4374; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4376 = 4'h9 == stack_num & 6'h3 == current_field_num ? field_stack_9_field_type_3_field_type :
    _GEN_4375; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4377 = 4'h9 == stack_num & 6'h4 == current_field_num ? field_stack_9_field_type_4_field_type :
    _GEN_4376; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4378 = 4'h9 == stack_num & 6'h5 == current_field_num ? field_stack_9_field_type_5_field_type :
    _GEN_4377; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4379 = 4'h9 == stack_num & 6'h6 == current_field_num ? field_stack_9_field_type_6_field_type :
    _GEN_4378; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4380 = 4'h9 == stack_num & 6'h7 == current_field_num ? field_stack_9_field_type_7_field_type :
    _GEN_4379; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4381 = 4'h9 == stack_num & 6'h8 == current_field_num ? field_stack_9_field_type_8_field_type :
    _GEN_4380; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4382 = 4'h9 == stack_num & 6'h9 == current_field_num ? field_stack_9_field_type_9_field_type :
    _GEN_4381; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4383 = 4'h9 == stack_num & 6'ha == current_field_num ? field_stack_9_field_type_10_field_type :
    _GEN_4382; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4384 = 4'h9 == stack_num & 6'hb == current_field_num ? field_stack_9_field_type_11_field_type :
    _GEN_4383; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4385 = 4'h9 == stack_num & 6'hc == current_field_num ? field_stack_9_field_type_12_field_type :
    _GEN_4384; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4386 = 4'h9 == stack_num & 6'hd == current_field_num ? field_stack_9_field_type_13_field_type :
    _GEN_4385; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4387 = 4'h9 == stack_num & 6'he == current_field_num ? field_stack_9_field_type_14_field_type :
    _GEN_4386; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4388 = 4'h9 == stack_num & 6'hf == current_field_num ? field_stack_9_field_type_15_field_type :
    _GEN_4387; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4389 = 4'h9 == stack_num & 6'h10 == current_field_num ? field_stack_9_field_type_16_field_type :
    _GEN_4388; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4390 = 4'h9 == stack_num & 6'h11 == current_field_num ? field_stack_9_field_type_17_field_type :
    _GEN_4389; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4391 = 4'h9 == stack_num & 6'h12 == current_field_num ? field_stack_9_field_type_18_field_type :
    _GEN_4390; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4392 = 4'h9 == stack_num & 6'h13 == current_field_num ? field_stack_9_field_type_19_field_type :
    _GEN_4391; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4393 = 4'h9 == stack_num & 6'h14 == current_field_num ? field_stack_9_field_type_20_field_type :
    _GEN_4392; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4394 = 4'h9 == stack_num & 6'h15 == current_field_num ? field_stack_9_field_type_21_field_type :
    _GEN_4393; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4395 = 4'h9 == stack_num & 6'h16 == current_field_num ? field_stack_9_field_type_22_field_type :
    _GEN_4394; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4396 = 4'h9 == stack_num & 6'h17 == current_field_num ? field_stack_9_field_type_23_field_type :
    _GEN_4395; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4397 = 4'h9 == stack_num & 6'h18 == current_field_num ? field_stack_9_field_type_24_field_type :
    _GEN_4396; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4398 = 4'h9 == stack_num & 6'h19 == current_field_num ? field_stack_9_field_type_25_field_type :
    _GEN_4397; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4399 = 4'h9 == stack_num & 6'h1a == current_field_num ? field_stack_9_field_type_26_field_type :
    _GEN_4398; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4400 = 4'h9 == stack_num & 6'h1b == current_field_num ? field_stack_9_field_type_27_field_type :
    _GEN_4399; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4401 = 4'h9 == stack_num & 6'h1c == current_field_num ? field_stack_9_field_type_28_field_type :
    _GEN_4400; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4402 = 4'h9 == stack_num & 6'h1d == current_field_num ? field_stack_9_field_type_29_field_type :
    _GEN_4401; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4403 = 4'h9 == stack_num & 6'h1e == current_field_num ? field_stack_9_field_type_30_field_type :
    _GEN_4402; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4404 = 4'h9 == stack_num & 6'h1f == current_field_num ? field_stack_9_field_type_31_field_type :
    _GEN_4403; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4405 = 4'h9 == stack_num & 6'h20 == current_field_num ? field_stack_9_field_type_32_field_type :
    _GEN_4404; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire  _GEN_11301 = 4'ha == stack_num; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4406 = 4'ha == stack_num & 6'h0 == current_field_num ? field_stack_10_field_type_0_field_type :
    _GEN_4405; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4407 = 4'ha == stack_num & 6'h1 == current_field_num ? field_stack_10_field_type_1_field_type :
    _GEN_4406; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4408 = 4'ha == stack_num & 6'h2 == current_field_num ? field_stack_10_field_type_2_field_type :
    _GEN_4407; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4409 = 4'ha == stack_num & 6'h3 == current_field_num ? field_stack_10_field_type_3_field_type :
    _GEN_4408; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4410 = 4'ha == stack_num & 6'h4 == current_field_num ? field_stack_10_field_type_4_field_type :
    _GEN_4409; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4411 = 4'ha == stack_num & 6'h5 == current_field_num ? field_stack_10_field_type_5_field_type :
    _GEN_4410; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4412 = 4'ha == stack_num & 6'h6 == current_field_num ? field_stack_10_field_type_6_field_type :
    _GEN_4411; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4413 = 4'ha == stack_num & 6'h7 == current_field_num ? field_stack_10_field_type_7_field_type :
    _GEN_4412; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4414 = 4'ha == stack_num & 6'h8 == current_field_num ? field_stack_10_field_type_8_field_type :
    _GEN_4413; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4415 = 4'ha == stack_num & 6'h9 == current_field_num ? field_stack_10_field_type_9_field_type :
    _GEN_4414; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4416 = 4'ha == stack_num & 6'ha == current_field_num ? field_stack_10_field_type_10_field_type :
    _GEN_4415; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4417 = 4'ha == stack_num & 6'hb == current_field_num ? field_stack_10_field_type_11_field_type :
    _GEN_4416; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4418 = 4'ha == stack_num & 6'hc == current_field_num ? field_stack_10_field_type_12_field_type :
    _GEN_4417; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4419 = 4'ha == stack_num & 6'hd == current_field_num ? field_stack_10_field_type_13_field_type :
    _GEN_4418; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4420 = 4'ha == stack_num & 6'he == current_field_num ? field_stack_10_field_type_14_field_type :
    _GEN_4419; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4421 = 4'ha == stack_num & 6'hf == current_field_num ? field_stack_10_field_type_15_field_type :
    _GEN_4420; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4422 = 4'ha == stack_num & 6'h10 == current_field_num ? field_stack_10_field_type_16_field_type :
    _GEN_4421; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4423 = 4'ha == stack_num & 6'h11 == current_field_num ? field_stack_10_field_type_17_field_type :
    _GEN_4422; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4424 = 4'ha == stack_num & 6'h12 == current_field_num ? field_stack_10_field_type_18_field_type :
    _GEN_4423; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4425 = 4'ha == stack_num & 6'h13 == current_field_num ? field_stack_10_field_type_19_field_type :
    _GEN_4424; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4426 = 4'ha == stack_num & 6'h14 == current_field_num ? field_stack_10_field_type_20_field_type :
    _GEN_4425; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4427 = 4'ha == stack_num & 6'h15 == current_field_num ? field_stack_10_field_type_21_field_type :
    _GEN_4426; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4428 = 4'ha == stack_num & 6'h16 == current_field_num ? field_stack_10_field_type_22_field_type :
    _GEN_4427; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4429 = 4'ha == stack_num & 6'h17 == current_field_num ? field_stack_10_field_type_23_field_type :
    _GEN_4428; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4430 = 4'ha == stack_num & 6'h18 == current_field_num ? field_stack_10_field_type_24_field_type :
    _GEN_4429; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4431 = 4'ha == stack_num & 6'h19 == current_field_num ? field_stack_10_field_type_25_field_type :
    _GEN_4430; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4432 = 4'ha == stack_num & 6'h1a == current_field_num ? field_stack_10_field_type_26_field_type :
    _GEN_4431; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4433 = 4'ha == stack_num & 6'h1b == current_field_num ? field_stack_10_field_type_27_field_type :
    _GEN_4432; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4434 = 4'ha == stack_num & 6'h1c == current_field_num ? field_stack_10_field_type_28_field_type :
    _GEN_4433; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4435 = 4'ha == stack_num & 6'h1d == current_field_num ? field_stack_10_field_type_29_field_type :
    _GEN_4434; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4436 = 4'ha == stack_num & 6'h1e == current_field_num ? field_stack_10_field_type_30_field_type :
    _GEN_4435; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4437 = 4'ha == stack_num & 6'h1f == current_field_num ? field_stack_10_field_type_31_field_type :
    _GEN_4436; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4438 = 4'ha == stack_num & 6'h20 == current_field_num ? field_stack_10_field_type_32_field_type :
    _GEN_4437; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire  _GEN_11367 = 4'hb == stack_num; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4439 = 4'hb == stack_num & 6'h0 == current_field_num ? field_stack_11_field_type_0_field_type :
    _GEN_4438; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4440 = 4'hb == stack_num & 6'h1 == current_field_num ? field_stack_11_field_type_1_field_type :
    _GEN_4439; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4441 = 4'hb == stack_num & 6'h2 == current_field_num ? field_stack_11_field_type_2_field_type :
    _GEN_4440; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4442 = 4'hb == stack_num & 6'h3 == current_field_num ? field_stack_11_field_type_3_field_type :
    _GEN_4441; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4443 = 4'hb == stack_num & 6'h4 == current_field_num ? field_stack_11_field_type_4_field_type :
    _GEN_4442; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4444 = 4'hb == stack_num & 6'h5 == current_field_num ? field_stack_11_field_type_5_field_type :
    _GEN_4443; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4445 = 4'hb == stack_num & 6'h6 == current_field_num ? field_stack_11_field_type_6_field_type :
    _GEN_4444; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4446 = 4'hb == stack_num & 6'h7 == current_field_num ? field_stack_11_field_type_7_field_type :
    _GEN_4445; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4447 = 4'hb == stack_num & 6'h8 == current_field_num ? field_stack_11_field_type_8_field_type :
    _GEN_4446; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4448 = 4'hb == stack_num & 6'h9 == current_field_num ? field_stack_11_field_type_9_field_type :
    _GEN_4447; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4449 = 4'hb == stack_num & 6'ha == current_field_num ? field_stack_11_field_type_10_field_type :
    _GEN_4448; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4450 = 4'hb == stack_num & 6'hb == current_field_num ? field_stack_11_field_type_11_field_type :
    _GEN_4449; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4451 = 4'hb == stack_num & 6'hc == current_field_num ? field_stack_11_field_type_12_field_type :
    _GEN_4450; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4452 = 4'hb == stack_num & 6'hd == current_field_num ? field_stack_11_field_type_13_field_type :
    _GEN_4451; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4453 = 4'hb == stack_num & 6'he == current_field_num ? field_stack_11_field_type_14_field_type :
    _GEN_4452; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4454 = 4'hb == stack_num & 6'hf == current_field_num ? field_stack_11_field_type_15_field_type :
    _GEN_4453; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4455 = 4'hb == stack_num & 6'h10 == current_field_num ? field_stack_11_field_type_16_field_type :
    _GEN_4454; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4456 = 4'hb == stack_num & 6'h11 == current_field_num ? field_stack_11_field_type_17_field_type :
    _GEN_4455; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4457 = 4'hb == stack_num & 6'h12 == current_field_num ? field_stack_11_field_type_18_field_type :
    _GEN_4456; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4458 = 4'hb == stack_num & 6'h13 == current_field_num ? field_stack_11_field_type_19_field_type :
    _GEN_4457; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4459 = 4'hb == stack_num & 6'h14 == current_field_num ? field_stack_11_field_type_20_field_type :
    _GEN_4458; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4460 = 4'hb == stack_num & 6'h15 == current_field_num ? field_stack_11_field_type_21_field_type :
    _GEN_4459; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4461 = 4'hb == stack_num & 6'h16 == current_field_num ? field_stack_11_field_type_22_field_type :
    _GEN_4460; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4462 = 4'hb == stack_num & 6'h17 == current_field_num ? field_stack_11_field_type_23_field_type :
    _GEN_4461; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4463 = 4'hb == stack_num & 6'h18 == current_field_num ? field_stack_11_field_type_24_field_type :
    _GEN_4462; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4464 = 4'hb == stack_num & 6'h19 == current_field_num ? field_stack_11_field_type_25_field_type :
    _GEN_4463; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4465 = 4'hb == stack_num & 6'h1a == current_field_num ? field_stack_11_field_type_26_field_type :
    _GEN_4464; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4466 = 4'hb == stack_num & 6'h1b == current_field_num ? field_stack_11_field_type_27_field_type :
    _GEN_4465; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4467 = 4'hb == stack_num & 6'h1c == current_field_num ? field_stack_11_field_type_28_field_type :
    _GEN_4466; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4468 = 4'hb == stack_num & 6'h1d == current_field_num ? field_stack_11_field_type_29_field_type :
    _GEN_4467; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4469 = 4'hb == stack_num & 6'h1e == current_field_num ? field_stack_11_field_type_30_field_type :
    _GEN_4468; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4470 = 4'hb == stack_num & 6'h1f == current_field_num ? field_stack_11_field_type_31_field_type :
    _GEN_4469; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4471 = 4'hb == stack_num & 6'h20 == current_field_num ? field_stack_11_field_type_32_field_type :
    _GEN_4470; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire  _GEN_11433 = 4'hc == stack_num; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4472 = 4'hc == stack_num & 6'h0 == current_field_num ? field_stack_12_field_type_0_field_type :
    _GEN_4471; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4473 = 4'hc == stack_num & 6'h1 == current_field_num ? field_stack_12_field_type_1_field_type :
    _GEN_4472; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4474 = 4'hc == stack_num & 6'h2 == current_field_num ? field_stack_12_field_type_2_field_type :
    _GEN_4473; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4475 = 4'hc == stack_num & 6'h3 == current_field_num ? field_stack_12_field_type_3_field_type :
    _GEN_4474; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4476 = 4'hc == stack_num & 6'h4 == current_field_num ? field_stack_12_field_type_4_field_type :
    _GEN_4475; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4477 = 4'hc == stack_num & 6'h5 == current_field_num ? field_stack_12_field_type_5_field_type :
    _GEN_4476; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4478 = 4'hc == stack_num & 6'h6 == current_field_num ? field_stack_12_field_type_6_field_type :
    _GEN_4477; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4479 = 4'hc == stack_num & 6'h7 == current_field_num ? field_stack_12_field_type_7_field_type :
    _GEN_4478; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4480 = 4'hc == stack_num & 6'h8 == current_field_num ? field_stack_12_field_type_8_field_type :
    _GEN_4479; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4481 = 4'hc == stack_num & 6'h9 == current_field_num ? field_stack_12_field_type_9_field_type :
    _GEN_4480; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4482 = 4'hc == stack_num & 6'ha == current_field_num ? field_stack_12_field_type_10_field_type :
    _GEN_4481; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4483 = 4'hc == stack_num & 6'hb == current_field_num ? field_stack_12_field_type_11_field_type :
    _GEN_4482; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4484 = 4'hc == stack_num & 6'hc == current_field_num ? field_stack_12_field_type_12_field_type :
    _GEN_4483; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4485 = 4'hc == stack_num & 6'hd == current_field_num ? field_stack_12_field_type_13_field_type :
    _GEN_4484; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4486 = 4'hc == stack_num & 6'he == current_field_num ? field_stack_12_field_type_14_field_type :
    _GEN_4485; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4487 = 4'hc == stack_num & 6'hf == current_field_num ? field_stack_12_field_type_15_field_type :
    _GEN_4486; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4488 = 4'hc == stack_num & 6'h10 == current_field_num ? field_stack_12_field_type_16_field_type :
    _GEN_4487; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4489 = 4'hc == stack_num & 6'h11 == current_field_num ? field_stack_12_field_type_17_field_type :
    _GEN_4488; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4490 = 4'hc == stack_num & 6'h12 == current_field_num ? field_stack_12_field_type_18_field_type :
    _GEN_4489; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4491 = 4'hc == stack_num & 6'h13 == current_field_num ? field_stack_12_field_type_19_field_type :
    _GEN_4490; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4492 = 4'hc == stack_num & 6'h14 == current_field_num ? field_stack_12_field_type_20_field_type :
    _GEN_4491; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4493 = 4'hc == stack_num & 6'h15 == current_field_num ? field_stack_12_field_type_21_field_type :
    _GEN_4492; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4494 = 4'hc == stack_num & 6'h16 == current_field_num ? field_stack_12_field_type_22_field_type :
    _GEN_4493; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4495 = 4'hc == stack_num & 6'h17 == current_field_num ? field_stack_12_field_type_23_field_type :
    _GEN_4494; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4496 = 4'hc == stack_num & 6'h18 == current_field_num ? field_stack_12_field_type_24_field_type :
    _GEN_4495; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4497 = 4'hc == stack_num & 6'h19 == current_field_num ? field_stack_12_field_type_25_field_type :
    _GEN_4496; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4498 = 4'hc == stack_num & 6'h1a == current_field_num ? field_stack_12_field_type_26_field_type :
    _GEN_4497; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4499 = 4'hc == stack_num & 6'h1b == current_field_num ? field_stack_12_field_type_27_field_type :
    _GEN_4498; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4500 = 4'hc == stack_num & 6'h1c == current_field_num ? field_stack_12_field_type_28_field_type :
    _GEN_4499; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4501 = 4'hc == stack_num & 6'h1d == current_field_num ? field_stack_12_field_type_29_field_type :
    _GEN_4500; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4502 = 4'hc == stack_num & 6'h1e == current_field_num ? field_stack_12_field_type_30_field_type :
    _GEN_4501; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4503 = 4'hc == stack_num & 6'h1f == current_field_num ? field_stack_12_field_type_31_field_type :
    _GEN_4502; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4504 = 4'hc == stack_num & 6'h20 == current_field_num ? field_stack_12_field_type_32_field_type :
    _GEN_4503; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire  _GEN_11499 = 4'hd == stack_num; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4505 = 4'hd == stack_num & 6'h0 == current_field_num ? field_stack_13_field_type_0_field_type :
    _GEN_4504; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4506 = 4'hd == stack_num & 6'h1 == current_field_num ? field_stack_13_field_type_1_field_type :
    _GEN_4505; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4507 = 4'hd == stack_num & 6'h2 == current_field_num ? field_stack_13_field_type_2_field_type :
    _GEN_4506; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4508 = 4'hd == stack_num & 6'h3 == current_field_num ? field_stack_13_field_type_3_field_type :
    _GEN_4507; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4509 = 4'hd == stack_num & 6'h4 == current_field_num ? field_stack_13_field_type_4_field_type :
    _GEN_4508; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4510 = 4'hd == stack_num & 6'h5 == current_field_num ? field_stack_13_field_type_5_field_type :
    _GEN_4509; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4511 = 4'hd == stack_num & 6'h6 == current_field_num ? field_stack_13_field_type_6_field_type :
    _GEN_4510; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4512 = 4'hd == stack_num & 6'h7 == current_field_num ? field_stack_13_field_type_7_field_type :
    _GEN_4511; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4513 = 4'hd == stack_num & 6'h8 == current_field_num ? field_stack_13_field_type_8_field_type :
    _GEN_4512; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4514 = 4'hd == stack_num & 6'h9 == current_field_num ? field_stack_13_field_type_9_field_type :
    _GEN_4513; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4515 = 4'hd == stack_num & 6'ha == current_field_num ? field_stack_13_field_type_10_field_type :
    _GEN_4514; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4516 = 4'hd == stack_num & 6'hb == current_field_num ? field_stack_13_field_type_11_field_type :
    _GEN_4515; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4517 = 4'hd == stack_num & 6'hc == current_field_num ? field_stack_13_field_type_12_field_type :
    _GEN_4516; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4518 = 4'hd == stack_num & 6'hd == current_field_num ? field_stack_13_field_type_13_field_type :
    _GEN_4517; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4519 = 4'hd == stack_num & 6'he == current_field_num ? field_stack_13_field_type_14_field_type :
    _GEN_4518; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4520 = 4'hd == stack_num & 6'hf == current_field_num ? field_stack_13_field_type_15_field_type :
    _GEN_4519; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4521 = 4'hd == stack_num & 6'h10 == current_field_num ? field_stack_13_field_type_16_field_type :
    _GEN_4520; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4522 = 4'hd == stack_num & 6'h11 == current_field_num ? field_stack_13_field_type_17_field_type :
    _GEN_4521; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4523 = 4'hd == stack_num & 6'h12 == current_field_num ? field_stack_13_field_type_18_field_type :
    _GEN_4522; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4524 = 4'hd == stack_num & 6'h13 == current_field_num ? field_stack_13_field_type_19_field_type :
    _GEN_4523; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4525 = 4'hd == stack_num & 6'h14 == current_field_num ? field_stack_13_field_type_20_field_type :
    _GEN_4524; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4526 = 4'hd == stack_num & 6'h15 == current_field_num ? field_stack_13_field_type_21_field_type :
    _GEN_4525; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4527 = 4'hd == stack_num & 6'h16 == current_field_num ? field_stack_13_field_type_22_field_type :
    _GEN_4526; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4528 = 4'hd == stack_num & 6'h17 == current_field_num ? field_stack_13_field_type_23_field_type :
    _GEN_4527; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4529 = 4'hd == stack_num & 6'h18 == current_field_num ? field_stack_13_field_type_24_field_type :
    _GEN_4528; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4530 = 4'hd == stack_num & 6'h19 == current_field_num ? field_stack_13_field_type_25_field_type :
    _GEN_4529; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4531 = 4'hd == stack_num & 6'h1a == current_field_num ? field_stack_13_field_type_26_field_type :
    _GEN_4530; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4532 = 4'hd == stack_num & 6'h1b == current_field_num ? field_stack_13_field_type_27_field_type :
    _GEN_4531; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4533 = 4'hd == stack_num & 6'h1c == current_field_num ? field_stack_13_field_type_28_field_type :
    _GEN_4532; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4534 = 4'hd == stack_num & 6'h1d == current_field_num ? field_stack_13_field_type_29_field_type :
    _GEN_4533; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4535 = 4'hd == stack_num & 6'h1e == current_field_num ? field_stack_13_field_type_30_field_type :
    _GEN_4534; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4536 = 4'hd == stack_num & 6'h1f == current_field_num ? field_stack_13_field_type_31_field_type :
    _GEN_4535; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4537 = 4'hd == stack_num & 6'h20 == current_field_num ? field_stack_13_field_type_32_field_type :
    _GEN_4536; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire  _GEN_11565 = 4'he == stack_num; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4538 = 4'he == stack_num & 6'h0 == current_field_num ? field_stack_14_field_type_0_field_type :
    _GEN_4537; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4539 = 4'he == stack_num & 6'h1 == current_field_num ? field_stack_14_field_type_1_field_type :
    _GEN_4538; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4540 = 4'he == stack_num & 6'h2 == current_field_num ? field_stack_14_field_type_2_field_type :
    _GEN_4539; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4541 = 4'he == stack_num & 6'h3 == current_field_num ? field_stack_14_field_type_3_field_type :
    _GEN_4540; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4542 = 4'he == stack_num & 6'h4 == current_field_num ? field_stack_14_field_type_4_field_type :
    _GEN_4541; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4543 = 4'he == stack_num & 6'h5 == current_field_num ? field_stack_14_field_type_5_field_type :
    _GEN_4542; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4544 = 4'he == stack_num & 6'h6 == current_field_num ? field_stack_14_field_type_6_field_type :
    _GEN_4543; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4545 = 4'he == stack_num & 6'h7 == current_field_num ? field_stack_14_field_type_7_field_type :
    _GEN_4544; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4546 = 4'he == stack_num & 6'h8 == current_field_num ? field_stack_14_field_type_8_field_type :
    _GEN_4545; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4547 = 4'he == stack_num & 6'h9 == current_field_num ? field_stack_14_field_type_9_field_type :
    _GEN_4546; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4548 = 4'he == stack_num & 6'ha == current_field_num ? field_stack_14_field_type_10_field_type :
    _GEN_4547; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4549 = 4'he == stack_num & 6'hb == current_field_num ? field_stack_14_field_type_11_field_type :
    _GEN_4548; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4550 = 4'he == stack_num & 6'hc == current_field_num ? field_stack_14_field_type_12_field_type :
    _GEN_4549; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4551 = 4'he == stack_num & 6'hd == current_field_num ? field_stack_14_field_type_13_field_type :
    _GEN_4550; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4552 = 4'he == stack_num & 6'he == current_field_num ? field_stack_14_field_type_14_field_type :
    _GEN_4551; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4553 = 4'he == stack_num & 6'hf == current_field_num ? field_stack_14_field_type_15_field_type :
    _GEN_4552; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4554 = 4'he == stack_num & 6'h10 == current_field_num ? field_stack_14_field_type_16_field_type :
    _GEN_4553; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4555 = 4'he == stack_num & 6'h11 == current_field_num ? field_stack_14_field_type_17_field_type :
    _GEN_4554; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4556 = 4'he == stack_num & 6'h12 == current_field_num ? field_stack_14_field_type_18_field_type :
    _GEN_4555; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4557 = 4'he == stack_num & 6'h13 == current_field_num ? field_stack_14_field_type_19_field_type :
    _GEN_4556; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4558 = 4'he == stack_num & 6'h14 == current_field_num ? field_stack_14_field_type_20_field_type :
    _GEN_4557; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4559 = 4'he == stack_num & 6'h15 == current_field_num ? field_stack_14_field_type_21_field_type :
    _GEN_4558; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4560 = 4'he == stack_num & 6'h16 == current_field_num ? field_stack_14_field_type_22_field_type :
    _GEN_4559; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4561 = 4'he == stack_num & 6'h17 == current_field_num ? field_stack_14_field_type_23_field_type :
    _GEN_4560; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4562 = 4'he == stack_num & 6'h18 == current_field_num ? field_stack_14_field_type_24_field_type :
    _GEN_4561; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4563 = 4'he == stack_num & 6'h19 == current_field_num ? field_stack_14_field_type_25_field_type :
    _GEN_4562; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4564 = 4'he == stack_num & 6'h1a == current_field_num ? field_stack_14_field_type_26_field_type :
    _GEN_4563; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4565 = 4'he == stack_num & 6'h1b == current_field_num ? field_stack_14_field_type_27_field_type :
    _GEN_4564; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4566 = 4'he == stack_num & 6'h1c == current_field_num ? field_stack_14_field_type_28_field_type :
    _GEN_4565; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4567 = 4'he == stack_num & 6'h1d == current_field_num ? field_stack_14_field_type_29_field_type :
    _GEN_4566; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4568 = 4'he == stack_num & 6'h1e == current_field_num ? field_stack_14_field_type_30_field_type :
    _GEN_4567; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4569 = 4'he == stack_num & 6'h1f == current_field_num ? field_stack_14_field_type_31_field_type :
    _GEN_4568; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [4:0] _GEN_4570 = 4'he == stack_num & 6'h20 == current_field_num ? field_stack_14_field_type_32_field_type :
    _GEN_4569; // @[Serializerhw.scala 136:89 Serializerhw.scala 136:89]
  wire [5:0] _current_field_num_T_1 = current_field_num - 6'h1; // @[Serializerhw.scala 138:66]
  wire [15:0] _GEN_5067 = _GEN_10643 & _GEN_10644 ? field_stack_0_field_type_1_sub_class_id :
    field_stack_0_field_type_0_sub_class_id; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5068 = _GEN_10643 & _GEN_10646 ? field_stack_0_field_type_2_sub_class_id : _GEN_5067; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5069 = _GEN_10643 & _GEN_10648 ? field_stack_0_field_type_3_sub_class_id : _GEN_5068; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5070 = _GEN_10643 & _GEN_10650 ? field_stack_0_field_type_4_sub_class_id : _GEN_5069; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5071 = _GEN_10643 & _GEN_10652 ? field_stack_0_field_type_5_sub_class_id : _GEN_5070; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5072 = _GEN_10643 & _GEN_10654 ? field_stack_0_field_type_6_sub_class_id : _GEN_5071; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5073 = _GEN_10643 & _GEN_10656 ? field_stack_0_field_type_7_sub_class_id : _GEN_5072; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5074 = _GEN_10643 & _GEN_10658 ? field_stack_0_field_type_8_sub_class_id : _GEN_5073; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5075 = _GEN_10643 & _GEN_10660 ? field_stack_0_field_type_9_sub_class_id : _GEN_5074; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5076 = _GEN_10643 & _GEN_10662 ? field_stack_0_field_type_10_sub_class_id : _GEN_5075; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5077 = _GEN_10643 & _GEN_10664 ? field_stack_0_field_type_11_sub_class_id : _GEN_5076; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5078 = _GEN_10643 & _GEN_10666 ? field_stack_0_field_type_12_sub_class_id : _GEN_5077; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5079 = _GEN_10643 & _GEN_10668 ? field_stack_0_field_type_13_sub_class_id : _GEN_5078; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5080 = _GEN_10643 & _GEN_10670 ? field_stack_0_field_type_14_sub_class_id : _GEN_5079; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5081 = _GEN_10643 & _GEN_10672 ? field_stack_0_field_type_15_sub_class_id : _GEN_5080; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5082 = _GEN_10643 & _GEN_10674 ? field_stack_0_field_type_16_sub_class_id : _GEN_5081; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5083 = _GEN_10643 & _GEN_10676 ? field_stack_0_field_type_17_sub_class_id : _GEN_5082; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5084 = _GEN_10643 & _GEN_10678 ? field_stack_0_field_type_18_sub_class_id : _GEN_5083; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5085 = _GEN_10643 & _GEN_10680 ? field_stack_0_field_type_19_sub_class_id : _GEN_5084; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5086 = _GEN_10643 & _GEN_10682 ? field_stack_0_field_type_20_sub_class_id : _GEN_5085; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5087 = _GEN_10643 & _GEN_10684 ? field_stack_0_field_type_21_sub_class_id : _GEN_5086; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5088 = _GEN_10643 & _GEN_10686 ? field_stack_0_field_type_22_sub_class_id : _GEN_5087; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5089 = _GEN_10643 & _GEN_10688 ? field_stack_0_field_type_23_sub_class_id : _GEN_5088; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5090 = _GEN_10643 & _GEN_10690 ? field_stack_0_field_type_24_sub_class_id : _GEN_5089; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5091 = _GEN_10643 & _GEN_10692 ? field_stack_0_field_type_25_sub_class_id : _GEN_5090; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5092 = _GEN_10643 & _GEN_10694 ? field_stack_0_field_type_26_sub_class_id : _GEN_5091; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5093 = _GEN_10643 & _GEN_10696 ? field_stack_0_field_type_27_sub_class_id : _GEN_5092; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5094 = _GEN_10643 & _GEN_10698 ? field_stack_0_field_type_28_sub_class_id : _GEN_5093; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5095 = _GEN_10643 & _GEN_10700 ? field_stack_0_field_type_29_sub_class_id : _GEN_5094; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5096 = _GEN_10643 & _GEN_10702 ? field_stack_0_field_type_30_sub_class_id : _GEN_5095; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5097 = _GEN_10643 & _GEN_10704 ? field_stack_0_field_type_31_sub_class_id : _GEN_5096; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5098 = _GEN_10643 & _GEN_10706 ? field_stack_0_field_type_32_sub_class_id : _GEN_5097; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5099 = _GEN_10707 & _GEN_10708 ? field_stack_1_field_type_0_sub_class_id : _GEN_5098; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5100 = _GEN_10707 & _GEN_10644 ? field_stack_1_field_type_1_sub_class_id : _GEN_5099; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5101 = _GEN_10707 & _GEN_10646 ? field_stack_1_field_type_2_sub_class_id : _GEN_5100; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5102 = _GEN_10707 & _GEN_10648 ? field_stack_1_field_type_3_sub_class_id : _GEN_5101; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5103 = _GEN_10707 & _GEN_10650 ? field_stack_1_field_type_4_sub_class_id : _GEN_5102; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5104 = _GEN_10707 & _GEN_10652 ? field_stack_1_field_type_5_sub_class_id : _GEN_5103; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5105 = _GEN_10707 & _GEN_10654 ? field_stack_1_field_type_6_sub_class_id : _GEN_5104; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5106 = _GEN_10707 & _GEN_10656 ? field_stack_1_field_type_7_sub_class_id : _GEN_5105; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5107 = _GEN_10707 & _GEN_10658 ? field_stack_1_field_type_8_sub_class_id : _GEN_5106; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5108 = _GEN_10707 & _GEN_10660 ? field_stack_1_field_type_9_sub_class_id : _GEN_5107; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5109 = _GEN_10707 & _GEN_10662 ? field_stack_1_field_type_10_sub_class_id : _GEN_5108; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5110 = _GEN_10707 & _GEN_10664 ? field_stack_1_field_type_11_sub_class_id : _GEN_5109; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5111 = _GEN_10707 & _GEN_10666 ? field_stack_1_field_type_12_sub_class_id : _GEN_5110; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5112 = _GEN_10707 & _GEN_10668 ? field_stack_1_field_type_13_sub_class_id : _GEN_5111; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5113 = _GEN_10707 & _GEN_10670 ? field_stack_1_field_type_14_sub_class_id : _GEN_5112; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5114 = _GEN_10707 & _GEN_10672 ? field_stack_1_field_type_15_sub_class_id : _GEN_5113; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5115 = _GEN_10707 & _GEN_10674 ? field_stack_1_field_type_16_sub_class_id : _GEN_5114; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5116 = _GEN_10707 & _GEN_10676 ? field_stack_1_field_type_17_sub_class_id : _GEN_5115; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5117 = _GEN_10707 & _GEN_10678 ? field_stack_1_field_type_18_sub_class_id : _GEN_5116; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5118 = _GEN_10707 & _GEN_10680 ? field_stack_1_field_type_19_sub_class_id : _GEN_5117; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5119 = _GEN_10707 & _GEN_10682 ? field_stack_1_field_type_20_sub_class_id : _GEN_5118; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5120 = _GEN_10707 & _GEN_10684 ? field_stack_1_field_type_21_sub_class_id : _GEN_5119; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5121 = _GEN_10707 & _GEN_10686 ? field_stack_1_field_type_22_sub_class_id : _GEN_5120; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5122 = _GEN_10707 & _GEN_10688 ? field_stack_1_field_type_23_sub_class_id : _GEN_5121; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5123 = _GEN_10707 & _GEN_10690 ? field_stack_1_field_type_24_sub_class_id : _GEN_5122; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5124 = _GEN_10707 & _GEN_10692 ? field_stack_1_field_type_25_sub_class_id : _GEN_5123; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5125 = _GEN_10707 & _GEN_10694 ? field_stack_1_field_type_26_sub_class_id : _GEN_5124; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5126 = _GEN_10707 & _GEN_10696 ? field_stack_1_field_type_27_sub_class_id : _GEN_5125; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5127 = _GEN_10707 & _GEN_10698 ? field_stack_1_field_type_28_sub_class_id : _GEN_5126; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5128 = _GEN_10707 & _GEN_10700 ? field_stack_1_field_type_29_sub_class_id : _GEN_5127; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5129 = _GEN_10707 & _GEN_10702 ? field_stack_1_field_type_30_sub_class_id : _GEN_5128; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5130 = _GEN_10707 & _GEN_10704 ? field_stack_1_field_type_31_sub_class_id : _GEN_5129; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5131 = _GEN_10707 & _GEN_10706 ? field_stack_1_field_type_32_sub_class_id : _GEN_5130; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5132 = _GEN_10773 & _GEN_10708 ? field_stack_2_field_type_0_sub_class_id : _GEN_5131; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5133 = _GEN_10773 & _GEN_10644 ? field_stack_2_field_type_1_sub_class_id : _GEN_5132; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5134 = _GEN_10773 & _GEN_10646 ? field_stack_2_field_type_2_sub_class_id : _GEN_5133; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5135 = _GEN_10773 & _GEN_10648 ? field_stack_2_field_type_3_sub_class_id : _GEN_5134; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5136 = _GEN_10773 & _GEN_10650 ? field_stack_2_field_type_4_sub_class_id : _GEN_5135; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5137 = _GEN_10773 & _GEN_10652 ? field_stack_2_field_type_5_sub_class_id : _GEN_5136; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5138 = _GEN_10773 & _GEN_10654 ? field_stack_2_field_type_6_sub_class_id : _GEN_5137; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5139 = _GEN_10773 & _GEN_10656 ? field_stack_2_field_type_7_sub_class_id : _GEN_5138; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5140 = _GEN_10773 & _GEN_10658 ? field_stack_2_field_type_8_sub_class_id : _GEN_5139; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5141 = _GEN_10773 & _GEN_10660 ? field_stack_2_field_type_9_sub_class_id : _GEN_5140; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5142 = _GEN_10773 & _GEN_10662 ? field_stack_2_field_type_10_sub_class_id : _GEN_5141; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5143 = _GEN_10773 & _GEN_10664 ? field_stack_2_field_type_11_sub_class_id : _GEN_5142; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5144 = _GEN_10773 & _GEN_10666 ? field_stack_2_field_type_12_sub_class_id : _GEN_5143; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5145 = _GEN_10773 & _GEN_10668 ? field_stack_2_field_type_13_sub_class_id : _GEN_5144; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5146 = _GEN_10773 & _GEN_10670 ? field_stack_2_field_type_14_sub_class_id : _GEN_5145; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5147 = _GEN_10773 & _GEN_10672 ? field_stack_2_field_type_15_sub_class_id : _GEN_5146; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5148 = _GEN_10773 & _GEN_10674 ? field_stack_2_field_type_16_sub_class_id : _GEN_5147; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5149 = _GEN_10773 & _GEN_10676 ? field_stack_2_field_type_17_sub_class_id : _GEN_5148; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5150 = _GEN_10773 & _GEN_10678 ? field_stack_2_field_type_18_sub_class_id : _GEN_5149; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5151 = _GEN_10773 & _GEN_10680 ? field_stack_2_field_type_19_sub_class_id : _GEN_5150; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5152 = _GEN_10773 & _GEN_10682 ? field_stack_2_field_type_20_sub_class_id : _GEN_5151; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5153 = _GEN_10773 & _GEN_10684 ? field_stack_2_field_type_21_sub_class_id : _GEN_5152; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5154 = _GEN_10773 & _GEN_10686 ? field_stack_2_field_type_22_sub_class_id : _GEN_5153; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5155 = _GEN_10773 & _GEN_10688 ? field_stack_2_field_type_23_sub_class_id : _GEN_5154; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5156 = _GEN_10773 & _GEN_10690 ? field_stack_2_field_type_24_sub_class_id : _GEN_5155; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5157 = _GEN_10773 & _GEN_10692 ? field_stack_2_field_type_25_sub_class_id : _GEN_5156; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5158 = _GEN_10773 & _GEN_10694 ? field_stack_2_field_type_26_sub_class_id : _GEN_5157; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5159 = _GEN_10773 & _GEN_10696 ? field_stack_2_field_type_27_sub_class_id : _GEN_5158; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5160 = _GEN_10773 & _GEN_10698 ? field_stack_2_field_type_28_sub_class_id : _GEN_5159; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5161 = _GEN_10773 & _GEN_10700 ? field_stack_2_field_type_29_sub_class_id : _GEN_5160; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5162 = _GEN_10773 & _GEN_10702 ? field_stack_2_field_type_30_sub_class_id : _GEN_5161; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5163 = _GEN_10773 & _GEN_10704 ? field_stack_2_field_type_31_sub_class_id : _GEN_5162; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5164 = _GEN_10773 & _GEN_10706 ? field_stack_2_field_type_32_sub_class_id : _GEN_5163; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5165 = _GEN_10839 & _GEN_10708 ? field_stack_3_field_type_0_sub_class_id : _GEN_5164; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5166 = _GEN_10839 & _GEN_10644 ? field_stack_3_field_type_1_sub_class_id : _GEN_5165; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5167 = _GEN_10839 & _GEN_10646 ? field_stack_3_field_type_2_sub_class_id : _GEN_5166; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5168 = _GEN_10839 & _GEN_10648 ? field_stack_3_field_type_3_sub_class_id : _GEN_5167; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5169 = _GEN_10839 & _GEN_10650 ? field_stack_3_field_type_4_sub_class_id : _GEN_5168; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5170 = _GEN_10839 & _GEN_10652 ? field_stack_3_field_type_5_sub_class_id : _GEN_5169; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5171 = _GEN_10839 & _GEN_10654 ? field_stack_3_field_type_6_sub_class_id : _GEN_5170; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5172 = _GEN_10839 & _GEN_10656 ? field_stack_3_field_type_7_sub_class_id : _GEN_5171; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5173 = _GEN_10839 & _GEN_10658 ? field_stack_3_field_type_8_sub_class_id : _GEN_5172; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5174 = _GEN_10839 & _GEN_10660 ? field_stack_3_field_type_9_sub_class_id : _GEN_5173; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5175 = _GEN_10839 & _GEN_10662 ? field_stack_3_field_type_10_sub_class_id : _GEN_5174; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5176 = _GEN_10839 & _GEN_10664 ? field_stack_3_field_type_11_sub_class_id : _GEN_5175; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5177 = _GEN_10839 & _GEN_10666 ? field_stack_3_field_type_12_sub_class_id : _GEN_5176; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5178 = _GEN_10839 & _GEN_10668 ? field_stack_3_field_type_13_sub_class_id : _GEN_5177; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5179 = _GEN_10839 & _GEN_10670 ? field_stack_3_field_type_14_sub_class_id : _GEN_5178; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5180 = _GEN_10839 & _GEN_10672 ? field_stack_3_field_type_15_sub_class_id : _GEN_5179; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5181 = _GEN_10839 & _GEN_10674 ? field_stack_3_field_type_16_sub_class_id : _GEN_5180; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5182 = _GEN_10839 & _GEN_10676 ? field_stack_3_field_type_17_sub_class_id : _GEN_5181; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5183 = _GEN_10839 & _GEN_10678 ? field_stack_3_field_type_18_sub_class_id : _GEN_5182; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5184 = _GEN_10839 & _GEN_10680 ? field_stack_3_field_type_19_sub_class_id : _GEN_5183; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5185 = _GEN_10839 & _GEN_10682 ? field_stack_3_field_type_20_sub_class_id : _GEN_5184; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5186 = _GEN_10839 & _GEN_10684 ? field_stack_3_field_type_21_sub_class_id : _GEN_5185; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5187 = _GEN_10839 & _GEN_10686 ? field_stack_3_field_type_22_sub_class_id : _GEN_5186; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5188 = _GEN_10839 & _GEN_10688 ? field_stack_3_field_type_23_sub_class_id : _GEN_5187; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5189 = _GEN_10839 & _GEN_10690 ? field_stack_3_field_type_24_sub_class_id : _GEN_5188; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5190 = _GEN_10839 & _GEN_10692 ? field_stack_3_field_type_25_sub_class_id : _GEN_5189; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5191 = _GEN_10839 & _GEN_10694 ? field_stack_3_field_type_26_sub_class_id : _GEN_5190; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5192 = _GEN_10839 & _GEN_10696 ? field_stack_3_field_type_27_sub_class_id : _GEN_5191; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5193 = _GEN_10839 & _GEN_10698 ? field_stack_3_field_type_28_sub_class_id : _GEN_5192; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5194 = _GEN_10839 & _GEN_10700 ? field_stack_3_field_type_29_sub_class_id : _GEN_5193; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5195 = _GEN_10839 & _GEN_10702 ? field_stack_3_field_type_30_sub_class_id : _GEN_5194; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5196 = _GEN_10839 & _GEN_10704 ? field_stack_3_field_type_31_sub_class_id : _GEN_5195; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5197 = _GEN_10839 & _GEN_10706 ? field_stack_3_field_type_32_sub_class_id : _GEN_5196; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5198 = _GEN_10905 & _GEN_10708 ? field_stack_4_field_type_0_sub_class_id : _GEN_5197; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5199 = _GEN_10905 & _GEN_10644 ? field_stack_4_field_type_1_sub_class_id : _GEN_5198; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5200 = _GEN_10905 & _GEN_10646 ? field_stack_4_field_type_2_sub_class_id : _GEN_5199; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5201 = _GEN_10905 & _GEN_10648 ? field_stack_4_field_type_3_sub_class_id : _GEN_5200; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5202 = _GEN_10905 & _GEN_10650 ? field_stack_4_field_type_4_sub_class_id : _GEN_5201; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5203 = _GEN_10905 & _GEN_10652 ? field_stack_4_field_type_5_sub_class_id : _GEN_5202; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5204 = _GEN_10905 & _GEN_10654 ? field_stack_4_field_type_6_sub_class_id : _GEN_5203; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5205 = _GEN_10905 & _GEN_10656 ? field_stack_4_field_type_7_sub_class_id : _GEN_5204; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5206 = _GEN_10905 & _GEN_10658 ? field_stack_4_field_type_8_sub_class_id : _GEN_5205; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5207 = _GEN_10905 & _GEN_10660 ? field_stack_4_field_type_9_sub_class_id : _GEN_5206; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5208 = _GEN_10905 & _GEN_10662 ? field_stack_4_field_type_10_sub_class_id : _GEN_5207; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5209 = _GEN_10905 & _GEN_10664 ? field_stack_4_field_type_11_sub_class_id : _GEN_5208; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5210 = _GEN_10905 & _GEN_10666 ? field_stack_4_field_type_12_sub_class_id : _GEN_5209; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5211 = _GEN_10905 & _GEN_10668 ? field_stack_4_field_type_13_sub_class_id : _GEN_5210; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5212 = _GEN_10905 & _GEN_10670 ? field_stack_4_field_type_14_sub_class_id : _GEN_5211; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5213 = _GEN_10905 & _GEN_10672 ? field_stack_4_field_type_15_sub_class_id : _GEN_5212; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5214 = _GEN_10905 & _GEN_10674 ? field_stack_4_field_type_16_sub_class_id : _GEN_5213; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5215 = _GEN_10905 & _GEN_10676 ? field_stack_4_field_type_17_sub_class_id : _GEN_5214; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5216 = _GEN_10905 & _GEN_10678 ? field_stack_4_field_type_18_sub_class_id : _GEN_5215; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5217 = _GEN_10905 & _GEN_10680 ? field_stack_4_field_type_19_sub_class_id : _GEN_5216; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5218 = _GEN_10905 & _GEN_10682 ? field_stack_4_field_type_20_sub_class_id : _GEN_5217; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5219 = _GEN_10905 & _GEN_10684 ? field_stack_4_field_type_21_sub_class_id : _GEN_5218; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5220 = _GEN_10905 & _GEN_10686 ? field_stack_4_field_type_22_sub_class_id : _GEN_5219; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5221 = _GEN_10905 & _GEN_10688 ? field_stack_4_field_type_23_sub_class_id : _GEN_5220; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5222 = _GEN_10905 & _GEN_10690 ? field_stack_4_field_type_24_sub_class_id : _GEN_5221; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5223 = _GEN_10905 & _GEN_10692 ? field_stack_4_field_type_25_sub_class_id : _GEN_5222; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5224 = _GEN_10905 & _GEN_10694 ? field_stack_4_field_type_26_sub_class_id : _GEN_5223; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5225 = _GEN_10905 & _GEN_10696 ? field_stack_4_field_type_27_sub_class_id : _GEN_5224; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5226 = _GEN_10905 & _GEN_10698 ? field_stack_4_field_type_28_sub_class_id : _GEN_5225; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5227 = _GEN_10905 & _GEN_10700 ? field_stack_4_field_type_29_sub_class_id : _GEN_5226; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5228 = _GEN_10905 & _GEN_10702 ? field_stack_4_field_type_30_sub_class_id : _GEN_5227; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5229 = _GEN_10905 & _GEN_10704 ? field_stack_4_field_type_31_sub_class_id : _GEN_5228; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5230 = _GEN_10905 & _GEN_10706 ? field_stack_4_field_type_32_sub_class_id : _GEN_5229; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5231 = _GEN_10971 & _GEN_10708 ? field_stack_5_field_type_0_sub_class_id : _GEN_5230; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5232 = _GEN_10971 & _GEN_10644 ? field_stack_5_field_type_1_sub_class_id : _GEN_5231; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5233 = _GEN_10971 & _GEN_10646 ? field_stack_5_field_type_2_sub_class_id : _GEN_5232; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5234 = _GEN_10971 & _GEN_10648 ? field_stack_5_field_type_3_sub_class_id : _GEN_5233; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5235 = _GEN_10971 & _GEN_10650 ? field_stack_5_field_type_4_sub_class_id : _GEN_5234; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5236 = _GEN_10971 & _GEN_10652 ? field_stack_5_field_type_5_sub_class_id : _GEN_5235; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5237 = _GEN_10971 & _GEN_10654 ? field_stack_5_field_type_6_sub_class_id : _GEN_5236; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5238 = _GEN_10971 & _GEN_10656 ? field_stack_5_field_type_7_sub_class_id : _GEN_5237; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5239 = _GEN_10971 & _GEN_10658 ? field_stack_5_field_type_8_sub_class_id : _GEN_5238; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5240 = _GEN_10971 & _GEN_10660 ? field_stack_5_field_type_9_sub_class_id : _GEN_5239; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5241 = _GEN_10971 & _GEN_10662 ? field_stack_5_field_type_10_sub_class_id : _GEN_5240; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5242 = _GEN_10971 & _GEN_10664 ? field_stack_5_field_type_11_sub_class_id : _GEN_5241; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5243 = _GEN_10971 & _GEN_10666 ? field_stack_5_field_type_12_sub_class_id : _GEN_5242; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5244 = _GEN_10971 & _GEN_10668 ? field_stack_5_field_type_13_sub_class_id : _GEN_5243; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5245 = _GEN_10971 & _GEN_10670 ? field_stack_5_field_type_14_sub_class_id : _GEN_5244; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5246 = _GEN_10971 & _GEN_10672 ? field_stack_5_field_type_15_sub_class_id : _GEN_5245; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5247 = _GEN_10971 & _GEN_10674 ? field_stack_5_field_type_16_sub_class_id : _GEN_5246; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5248 = _GEN_10971 & _GEN_10676 ? field_stack_5_field_type_17_sub_class_id : _GEN_5247; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5249 = _GEN_10971 & _GEN_10678 ? field_stack_5_field_type_18_sub_class_id : _GEN_5248; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5250 = _GEN_10971 & _GEN_10680 ? field_stack_5_field_type_19_sub_class_id : _GEN_5249; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5251 = _GEN_10971 & _GEN_10682 ? field_stack_5_field_type_20_sub_class_id : _GEN_5250; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5252 = _GEN_10971 & _GEN_10684 ? field_stack_5_field_type_21_sub_class_id : _GEN_5251; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5253 = _GEN_10971 & _GEN_10686 ? field_stack_5_field_type_22_sub_class_id : _GEN_5252; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5254 = _GEN_10971 & _GEN_10688 ? field_stack_5_field_type_23_sub_class_id : _GEN_5253; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5255 = _GEN_10971 & _GEN_10690 ? field_stack_5_field_type_24_sub_class_id : _GEN_5254; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5256 = _GEN_10971 & _GEN_10692 ? field_stack_5_field_type_25_sub_class_id : _GEN_5255; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5257 = _GEN_10971 & _GEN_10694 ? field_stack_5_field_type_26_sub_class_id : _GEN_5256; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5258 = _GEN_10971 & _GEN_10696 ? field_stack_5_field_type_27_sub_class_id : _GEN_5257; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5259 = _GEN_10971 & _GEN_10698 ? field_stack_5_field_type_28_sub_class_id : _GEN_5258; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5260 = _GEN_10971 & _GEN_10700 ? field_stack_5_field_type_29_sub_class_id : _GEN_5259; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5261 = _GEN_10971 & _GEN_10702 ? field_stack_5_field_type_30_sub_class_id : _GEN_5260; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5262 = _GEN_10971 & _GEN_10704 ? field_stack_5_field_type_31_sub_class_id : _GEN_5261; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5263 = _GEN_10971 & _GEN_10706 ? field_stack_5_field_type_32_sub_class_id : _GEN_5262; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5264 = _GEN_11037 & _GEN_10708 ? field_stack_6_field_type_0_sub_class_id : _GEN_5263; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5265 = _GEN_11037 & _GEN_10644 ? field_stack_6_field_type_1_sub_class_id : _GEN_5264; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5266 = _GEN_11037 & _GEN_10646 ? field_stack_6_field_type_2_sub_class_id : _GEN_5265; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5267 = _GEN_11037 & _GEN_10648 ? field_stack_6_field_type_3_sub_class_id : _GEN_5266; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5268 = _GEN_11037 & _GEN_10650 ? field_stack_6_field_type_4_sub_class_id : _GEN_5267; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5269 = _GEN_11037 & _GEN_10652 ? field_stack_6_field_type_5_sub_class_id : _GEN_5268; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5270 = _GEN_11037 & _GEN_10654 ? field_stack_6_field_type_6_sub_class_id : _GEN_5269; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5271 = _GEN_11037 & _GEN_10656 ? field_stack_6_field_type_7_sub_class_id : _GEN_5270; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5272 = _GEN_11037 & _GEN_10658 ? field_stack_6_field_type_8_sub_class_id : _GEN_5271; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5273 = _GEN_11037 & _GEN_10660 ? field_stack_6_field_type_9_sub_class_id : _GEN_5272; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5274 = _GEN_11037 & _GEN_10662 ? field_stack_6_field_type_10_sub_class_id : _GEN_5273; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5275 = _GEN_11037 & _GEN_10664 ? field_stack_6_field_type_11_sub_class_id : _GEN_5274; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5276 = _GEN_11037 & _GEN_10666 ? field_stack_6_field_type_12_sub_class_id : _GEN_5275; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5277 = _GEN_11037 & _GEN_10668 ? field_stack_6_field_type_13_sub_class_id : _GEN_5276; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5278 = _GEN_11037 & _GEN_10670 ? field_stack_6_field_type_14_sub_class_id : _GEN_5277; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5279 = _GEN_11037 & _GEN_10672 ? field_stack_6_field_type_15_sub_class_id : _GEN_5278; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5280 = _GEN_11037 & _GEN_10674 ? field_stack_6_field_type_16_sub_class_id : _GEN_5279; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5281 = _GEN_11037 & _GEN_10676 ? field_stack_6_field_type_17_sub_class_id : _GEN_5280; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5282 = _GEN_11037 & _GEN_10678 ? field_stack_6_field_type_18_sub_class_id : _GEN_5281; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5283 = _GEN_11037 & _GEN_10680 ? field_stack_6_field_type_19_sub_class_id : _GEN_5282; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5284 = _GEN_11037 & _GEN_10682 ? field_stack_6_field_type_20_sub_class_id : _GEN_5283; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5285 = _GEN_11037 & _GEN_10684 ? field_stack_6_field_type_21_sub_class_id : _GEN_5284; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5286 = _GEN_11037 & _GEN_10686 ? field_stack_6_field_type_22_sub_class_id : _GEN_5285; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5287 = _GEN_11037 & _GEN_10688 ? field_stack_6_field_type_23_sub_class_id : _GEN_5286; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5288 = _GEN_11037 & _GEN_10690 ? field_stack_6_field_type_24_sub_class_id : _GEN_5287; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5289 = _GEN_11037 & _GEN_10692 ? field_stack_6_field_type_25_sub_class_id : _GEN_5288; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5290 = _GEN_11037 & _GEN_10694 ? field_stack_6_field_type_26_sub_class_id : _GEN_5289; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5291 = _GEN_11037 & _GEN_10696 ? field_stack_6_field_type_27_sub_class_id : _GEN_5290; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5292 = _GEN_11037 & _GEN_10698 ? field_stack_6_field_type_28_sub_class_id : _GEN_5291; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5293 = _GEN_11037 & _GEN_10700 ? field_stack_6_field_type_29_sub_class_id : _GEN_5292; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5294 = _GEN_11037 & _GEN_10702 ? field_stack_6_field_type_30_sub_class_id : _GEN_5293; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5295 = _GEN_11037 & _GEN_10704 ? field_stack_6_field_type_31_sub_class_id : _GEN_5294; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5296 = _GEN_11037 & _GEN_10706 ? field_stack_6_field_type_32_sub_class_id : _GEN_5295; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5297 = _GEN_11103 & _GEN_10708 ? field_stack_7_field_type_0_sub_class_id : _GEN_5296; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5298 = _GEN_11103 & _GEN_10644 ? field_stack_7_field_type_1_sub_class_id : _GEN_5297; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5299 = _GEN_11103 & _GEN_10646 ? field_stack_7_field_type_2_sub_class_id : _GEN_5298; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5300 = _GEN_11103 & _GEN_10648 ? field_stack_7_field_type_3_sub_class_id : _GEN_5299; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5301 = _GEN_11103 & _GEN_10650 ? field_stack_7_field_type_4_sub_class_id : _GEN_5300; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5302 = _GEN_11103 & _GEN_10652 ? field_stack_7_field_type_5_sub_class_id : _GEN_5301; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5303 = _GEN_11103 & _GEN_10654 ? field_stack_7_field_type_6_sub_class_id : _GEN_5302; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5304 = _GEN_11103 & _GEN_10656 ? field_stack_7_field_type_7_sub_class_id : _GEN_5303; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5305 = _GEN_11103 & _GEN_10658 ? field_stack_7_field_type_8_sub_class_id : _GEN_5304; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5306 = _GEN_11103 & _GEN_10660 ? field_stack_7_field_type_9_sub_class_id : _GEN_5305; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5307 = _GEN_11103 & _GEN_10662 ? field_stack_7_field_type_10_sub_class_id : _GEN_5306; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5308 = _GEN_11103 & _GEN_10664 ? field_stack_7_field_type_11_sub_class_id : _GEN_5307; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5309 = _GEN_11103 & _GEN_10666 ? field_stack_7_field_type_12_sub_class_id : _GEN_5308; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5310 = _GEN_11103 & _GEN_10668 ? field_stack_7_field_type_13_sub_class_id : _GEN_5309; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5311 = _GEN_11103 & _GEN_10670 ? field_stack_7_field_type_14_sub_class_id : _GEN_5310; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5312 = _GEN_11103 & _GEN_10672 ? field_stack_7_field_type_15_sub_class_id : _GEN_5311; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5313 = _GEN_11103 & _GEN_10674 ? field_stack_7_field_type_16_sub_class_id : _GEN_5312; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5314 = _GEN_11103 & _GEN_10676 ? field_stack_7_field_type_17_sub_class_id : _GEN_5313; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5315 = _GEN_11103 & _GEN_10678 ? field_stack_7_field_type_18_sub_class_id : _GEN_5314; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5316 = _GEN_11103 & _GEN_10680 ? field_stack_7_field_type_19_sub_class_id : _GEN_5315; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5317 = _GEN_11103 & _GEN_10682 ? field_stack_7_field_type_20_sub_class_id : _GEN_5316; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5318 = _GEN_11103 & _GEN_10684 ? field_stack_7_field_type_21_sub_class_id : _GEN_5317; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5319 = _GEN_11103 & _GEN_10686 ? field_stack_7_field_type_22_sub_class_id : _GEN_5318; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5320 = _GEN_11103 & _GEN_10688 ? field_stack_7_field_type_23_sub_class_id : _GEN_5319; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5321 = _GEN_11103 & _GEN_10690 ? field_stack_7_field_type_24_sub_class_id : _GEN_5320; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5322 = _GEN_11103 & _GEN_10692 ? field_stack_7_field_type_25_sub_class_id : _GEN_5321; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5323 = _GEN_11103 & _GEN_10694 ? field_stack_7_field_type_26_sub_class_id : _GEN_5322; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5324 = _GEN_11103 & _GEN_10696 ? field_stack_7_field_type_27_sub_class_id : _GEN_5323; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5325 = _GEN_11103 & _GEN_10698 ? field_stack_7_field_type_28_sub_class_id : _GEN_5324; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5326 = _GEN_11103 & _GEN_10700 ? field_stack_7_field_type_29_sub_class_id : _GEN_5325; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5327 = _GEN_11103 & _GEN_10702 ? field_stack_7_field_type_30_sub_class_id : _GEN_5326; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5328 = _GEN_11103 & _GEN_10704 ? field_stack_7_field_type_31_sub_class_id : _GEN_5327; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5329 = _GEN_11103 & _GEN_10706 ? field_stack_7_field_type_32_sub_class_id : _GEN_5328; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5330 = _GEN_11169 & _GEN_10708 ? field_stack_8_field_type_0_sub_class_id : _GEN_5329; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5331 = _GEN_11169 & _GEN_10644 ? field_stack_8_field_type_1_sub_class_id : _GEN_5330; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5332 = _GEN_11169 & _GEN_10646 ? field_stack_8_field_type_2_sub_class_id : _GEN_5331; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5333 = _GEN_11169 & _GEN_10648 ? field_stack_8_field_type_3_sub_class_id : _GEN_5332; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5334 = _GEN_11169 & _GEN_10650 ? field_stack_8_field_type_4_sub_class_id : _GEN_5333; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5335 = _GEN_11169 & _GEN_10652 ? field_stack_8_field_type_5_sub_class_id : _GEN_5334; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5336 = _GEN_11169 & _GEN_10654 ? field_stack_8_field_type_6_sub_class_id : _GEN_5335; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5337 = _GEN_11169 & _GEN_10656 ? field_stack_8_field_type_7_sub_class_id : _GEN_5336; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5338 = _GEN_11169 & _GEN_10658 ? field_stack_8_field_type_8_sub_class_id : _GEN_5337; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5339 = _GEN_11169 & _GEN_10660 ? field_stack_8_field_type_9_sub_class_id : _GEN_5338; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5340 = _GEN_11169 & _GEN_10662 ? field_stack_8_field_type_10_sub_class_id : _GEN_5339; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5341 = _GEN_11169 & _GEN_10664 ? field_stack_8_field_type_11_sub_class_id : _GEN_5340; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5342 = _GEN_11169 & _GEN_10666 ? field_stack_8_field_type_12_sub_class_id : _GEN_5341; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5343 = _GEN_11169 & _GEN_10668 ? field_stack_8_field_type_13_sub_class_id : _GEN_5342; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5344 = _GEN_11169 & _GEN_10670 ? field_stack_8_field_type_14_sub_class_id : _GEN_5343; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5345 = _GEN_11169 & _GEN_10672 ? field_stack_8_field_type_15_sub_class_id : _GEN_5344; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5346 = _GEN_11169 & _GEN_10674 ? field_stack_8_field_type_16_sub_class_id : _GEN_5345; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5347 = _GEN_11169 & _GEN_10676 ? field_stack_8_field_type_17_sub_class_id : _GEN_5346; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5348 = _GEN_11169 & _GEN_10678 ? field_stack_8_field_type_18_sub_class_id : _GEN_5347; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5349 = _GEN_11169 & _GEN_10680 ? field_stack_8_field_type_19_sub_class_id : _GEN_5348; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5350 = _GEN_11169 & _GEN_10682 ? field_stack_8_field_type_20_sub_class_id : _GEN_5349; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5351 = _GEN_11169 & _GEN_10684 ? field_stack_8_field_type_21_sub_class_id : _GEN_5350; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5352 = _GEN_11169 & _GEN_10686 ? field_stack_8_field_type_22_sub_class_id : _GEN_5351; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5353 = _GEN_11169 & _GEN_10688 ? field_stack_8_field_type_23_sub_class_id : _GEN_5352; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5354 = _GEN_11169 & _GEN_10690 ? field_stack_8_field_type_24_sub_class_id : _GEN_5353; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5355 = _GEN_11169 & _GEN_10692 ? field_stack_8_field_type_25_sub_class_id : _GEN_5354; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5356 = _GEN_11169 & _GEN_10694 ? field_stack_8_field_type_26_sub_class_id : _GEN_5355; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5357 = _GEN_11169 & _GEN_10696 ? field_stack_8_field_type_27_sub_class_id : _GEN_5356; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5358 = _GEN_11169 & _GEN_10698 ? field_stack_8_field_type_28_sub_class_id : _GEN_5357; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5359 = _GEN_11169 & _GEN_10700 ? field_stack_8_field_type_29_sub_class_id : _GEN_5358; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5360 = _GEN_11169 & _GEN_10702 ? field_stack_8_field_type_30_sub_class_id : _GEN_5359; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5361 = _GEN_11169 & _GEN_10704 ? field_stack_8_field_type_31_sub_class_id : _GEN_5360; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5362 = _GEN_11169 & _GEN_10706 ? field_stack_8_field_type_32_sub_class_id : _GEN_5361; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5363 = _GEN_11235 & _GEN_10708 ? field_stack_9_field_type_0_sub_class_id : _GEN_5362; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5364 = _GEN_11235 & _GEN_10644 ? field_stack_9_field_type_1_sub_class_id : _GEN_5363; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5365 = _GEN_11235 & _GEN_10646 ? field_stack_9_field_type_2_sub_class_id : _GEN_5364; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5366 = _GEN_11235 & _GEN_10648 ? field_stack_9_field_type_3_sub_class_id : _GEN_5365; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5367 = _GEN_11235 & _GEN_10650 ? field_stack_9_field_type_4_sub_class_id : _GEN_5366; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5368 = _GEN_11235 & _GEN_10652 ? field_stack_9_field_type_5_sub_class_id : _GEN_5367; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5369 = _GEN_11235 & _GEN_10654 ? field_stack_9_field_type_6_sub_class_id : _GEN_5368; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5370 = _GEN_11235 & _GEN_10656 ? field_stack_9_field_type_7_sub_class_id : _GEN_5369; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5371 = _GEN_11235 & _GEN_10658 ? field_stack_9_field_type_8_sub_class_id : _GEN_5370; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5372 = _GEN_11235 & _GEN_10660 ? field_stack_9_field_type_9_sub_class_id : _GEN_5371; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5373 = _GEN_11235 & _GEN_10662 ? field_stack_9_field_type_10_sub_class_id : _GEN_5372; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5374 = _GEN_11235 & _GEN_10664 ? field_stack_9_field_type_11_sub_class_id : _GEN_5373; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5375 = _GEN_11235 & _GEN_10666 ? field_stack_9_field_type_12_sub_class_id : _GEN_5374; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5376 = _GEN_11235 & _GEN_10668 ? field_stack_9_field_type_13_sub_class_id : _GEN_5375; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5377 = _GEN_11235 & _GEN_10670 ? field_stack_9_field_type_14_sub_class_id : _GEN_5376; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5378 = _GEN_11235 & _GEN_10672 ? field_stack_9_field_type_15_sub_class_id : _GEN_5377; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5379 = _GEN_11235 & _GEN_10674 ? field_stack_9_field_type_16_sub_class_id : _GEN_5378; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5380 = _GEN_11235 & _GEN_10676 ? field_stack_9_field_type_17_sub_class_id : _GEN_5379; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5381 = _GEN_11235 & _GEN_10678 ? field_stack_9_field_type_18_sub_class_id : _GEN_5380; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5382 = _GEN_11235 & _GEN_10680 ? field_stack_9_field_type_19_sub_class_id : _GEN_5381; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5383 = _GEN_11235 & _GEN_10682 ? field_stack_9_field_type_20_sub_class_id : _GEN_5382; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5384 = _GEN_11235 & _GEN_10684 ? field_stack_9_field_type_21_sub_class_id : _GEN_5383; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5385 = _GEN_11235 & _GEN_10686 ? field_stack_9_field_type_22_sub_class_id : _GEN_5384; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5386 = _GEN_11235 & _GEN_10688 ? field_stack_9_field_type_23_sub_class_id : _GEN_5385; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5387 = _GEN_11235 & _GEN_10690 ? field_stack_9_field_type_24_sub_class_id : _GEN_5386; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5388 = _GEN_11235 & _GEN_10692 ? field_stack_9_field_type_25_sub_class_id : _GEN_5387; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5389 = _GEN_11235 & _GEN_10694 ? field_stack_9_field_type_26_sub_class_id : _GEN_5388; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5390 = _GEN_11235 & _GEN_10696 ? field_stack_9_field_type_27_sub_class_id : _GEN_5389; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5391 = _GEN_11235 & _GEN_10698 ? field_stack_9_field_type_28_sub_class_id : _GEN_5390; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5392 = _GEN_11235 & _GEN_10700 ? field_stack_9_field_type_29_sub_class_id : _GEN_5391; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5393 = _GEN_11235 & _GEN_10702 ? field_stack_9_field_type_30_sub_class_id : _GEN_5392; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5394 = _GEN_11235 & _GEN_10704 ? field_stack_9_field_type_31_sub_class_id : _GEN_5393; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5395 = _GEN_11235 & _GEN_10706 ? field_stack_9_field_type_32_sub_class_id : _GEN_5394; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5396 = _GEN_11301 & _GEN_10708 ? field_stack_10_field_type_0_sub_class_id : _GEN_5395; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5397 = _GEN_11301 & _GEN_10644 ? field_stack_10_field_type_1_sub_class_id : _GEN_5396; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5398 = _GEN_11301 & _GEN_10646 ? field_stack_10_field_type_2_sub_class_id : _GEN_5397; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5399 = _GEN_11301 & _GEN_10648 ? field_stack_10_field_type_3_sub_class_id : _GEN_5398; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5400 = _GEN_11301 & _GEN_10650 ? field_stack_10_field_type_4_sub_class_id : _GEN_5399; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5401 = _GEN_11301 & _GEN_10652 ? field_stack_10_field_type_5_sub_class_id : _GEN_5400; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5402 = _GEN_11301 & _GEN_10654 ? field_stack_10_field_type_6_sub_class_id : _GEN_5401; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5403 = _GEN_11301 & _GEN_10656 ? field_stack_10_field_type_7_sub_class_id : _GEN_5402; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5404 = _GEN_11301 & _GEN_10658 ? field_stack_10_field_type_8_sub_class_id : _GEN_5403; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5405 = _GEN_11301 & _GEN_10660 ? field_stack_10_field_type_9_sub_class_id : _GEN_5404; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5406 = _GEN_11301 & _GEN_10662 ? field_stack_10_field_type_10_sub_class_id : _GEN_5405; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5407 = _GEN_11301 & _GEN_10664 ? field_stack_10_field_type_11_sub_class_id : _GEN_5406; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5408 = _GEN_11301 & _GEN_10666 ? field_stack_10_field_type_12_sub_class_id : _GEN_5407; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5409 = _GEN_11301 & _GEN_10668 ? field_stack_10_field_type_13_sub_class_id : _GEN_5408; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5410 = _GEN_11301 & _GEN_10670 ? field_stack_10_field_type_14_sub_class_id : _GEN_5409; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5411 = _GEN_11301 & _GEN_10672 ? field_stack_10_field_type_15_sub_class_id : _GEN_5410; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5412 = _GEN_11301 & _GEN_10674 ? field_stack_10_field_type_16_sub_class_id : _GEN_5411; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5413 = _GEN_11301 & _GEN_10676 ? field_stack_10_field_type_17_sub_class_id : _GEN_5412; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5414 = _GEN_11301 & _GEN_10678 ? field_stack_10_field_type_18_sub_class_id : _GEN_5413; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5415 = _GEN_11301 & _GEN_10680 ? field_stack_10_field_type_19_sub_class_id : _GEN_5414; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5416 = _GEN_11301 & _GEN_10682 ? field_stack_10_field_type_20_sub_class_id : _GEN_5415; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5417 = _GEN_11301 & _GEN_10684 ? field_stack_10_field_type_21_sub_class_id : _GEN_5416; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5418 = _GEN_11301 & _GEN_10686 ? field_stack_10_field_type_22_sub_class_id : _GEN_5417; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5419 = _GEN_11301 & _GEN_10688 ? field_stack_10_field_type_23_sub_class_id : _GEN_5418; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5420 = _GEN_11301 & _GEN_10690 ? field_stack_10_field_type_24_sub_class_id : _GEN_5419; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5421 = _GEN_11301 & _GEN_10692 ? field_stack_10_field_type_25_sub_class_id : _GEN_5420; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5422 = _GEN_11301 & _GEN_10694 ? field_stack_10_field_type_26_sub_class_id : _GEN_5421; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5423 = _GEN_11301 & _GEN_10696 ? field_stack_10_field_type_27_sub_class_id : _GEN_5422; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5424 = _GEN_11301 & _GEN_10698 ? field_stack_10_field_type_28_sub_class_id : _GEN_5423; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5425 = _GEN_11301 & _GEN_10700 ? field_stack_10_field_type_29_sub_class_id : _GEN_5424; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5426 = _GEN_11301 & _GEN_10702 ? field_stack_10_field_type_30_sub_class_id : _GEN_5425; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5427 = _GEN_11301 & _GEN_10704 ? field_stack_10_field_type_31_sub_class_id : _GEN_5426; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5428 = _GEN_11301 & _GEN_10706 ? field_stack_10_field_type_32_sub_class_id : _GEN_5427; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5429 = _GEN_11367 & _GEN_10708 ? field_stack_11_field_type_0_sub_class_id : _GEN_5428; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5430 = _GEN_11367 & _GEN_10644 ? field_stack_11_field_type_1_sub_class_id : _GEN_5429; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5431 = _GEN_11367 & _GEN_10646 ? field_stack_11_field_type_2_sub_class_id : _GEN_5430; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5432 = _GEN_11367 & _GEN_10648 ? field_stack_11_field_type_3_sub_class_id : _GEN_5431; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5433 = _GEN_11367 & _GEN_10650 ? field_stack_11_field_type_4_sub_class_id : _GEN_5432; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5434 = _GEN_11367 & _GEN_10652 ? field_stack_11_field_type_5_sub_class_id : _GEN_5433; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5435 = _GEN_11367 & _GEN_10654 ? field_stack_11_field_type_6_sub_class_id : _GEN_5434; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5436 = _GEN_11367 & _GEN_10656 ? field_stack_11_field_type_7_sub_class_id : _GEN_5435; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5437 = _GEN_11367 & _GEN_10658 ? field_stack_11_field_type_8_sub_class_id : _GEN_5436; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5438 = _GEN_11367 & _GEN_10660 ? field_stack_11_field_type_9_sub_class_id : _GEN_5437; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5439 = _GEN_11367 & _GEN_10662 ? field_stack_11_field_type_10_sub_class_id : _GEN_5438; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5440 = _GEN_11367 & _GEN_10664 ? field_stack_11_field_type_11_sub_class_id : _GEN_5439; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5441 = _GEN_11367 & _GEN_10666 ? field_stack_11_field_type_12_sub_class_id : _GEN_5440; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5442 = _GEN_11367 & _GEN_10668 ? field_stack_11_field_type_13_sub_class_id : _GEN_5441; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5443 = _GEN_11367 & _GEN_10670 ? field_stack_11_field_type_14_sub_class_id : _GEN_5442; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5444 = _GEN_11367 & _GEN_10672 ? field_stack_11_field_type_15_sub_class_id : _GEN_5443; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5445 = _GEN_11367 & _GEN_10674 ? field_stack_11_field_type_16_sub_class_id : _GEN_5444; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5446 = _GEN_11367 & _GEN_10676 ? field_stack_11_field_type_17_sub_class_id : _GEN_5445; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5447 = _GEN_11367 & _GEN_10678 ? field_stack_11_field_type_18_sub_class_id : _GEN_5446; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5448 = _GEN_11367 & _GEN_10680 ? field_stack_11_field_type_19_sub_class_id : _GEN_5447; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5449 = _GEN_11367 & _GEN_10682 ? field_stack_11_field_type_20_sub_class_id : _GEN_5448; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5450 = _GEN_11367 & _GEN_10684 ? field_stack_11_field_type_21_sub_class_id : _GEN_5449; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5451 = _GEN_11367 & _GEN_10686 ? field_stack_11_field_type_22_sub_class_id : _GEN_5450; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5452 = _GEN_11367 & _GEN_10688 ? field_stack_11_field_type_23_sub_class_id : _GEN_5451; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5453 = _GEN_11367 & _GEN_10690 ? field_stack_11_field_type_24_sub_class_id : _GEN_5452; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5454 = _GEN_11367 & _GEN_10692 ? field_stack_11_field_type_25_sub_class_id : _GEN_5453; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5455 = _GEN_11367 & _GEN_10694 ? field_stack_11_field_type_26_sub_class_id : _GEN_5454; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5456 = _GEN_11367 & _GEN_10696 ? field_stack_11_field_type_27_sub_class_id : _GEN_5455; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5457 = _GEN_11367 & _GEN_10698 ? field_stack_11_field_type_28_sub_class_id : _GEN_5456; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5458 = _GEN_11367 & _GEN_10700 ? field_stack_11_field_type_29_sub_class_id : _GEN_5457; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5459 = _GEN_11367 & _GEN_10702 ? field_stack_11_field_type_30_sub_class_id : _GEN_5458; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5460 = _GEN_11367 & _GEN_10704 ? field_stack_11_field_type_31_sub_class_id : _GEN_5459; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5461 = _GEN_11367 & _GEN_10706 ? field_stack_11_field_type_32_sub_class_id : _GEN_5460; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5462 = _GEN_11433 & _GEN_10708 ? field_stack_12_field_type_0_sub_class_id : _GEN_5461; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5463 = _GEN_11433 & _GEN_10644 ? field_stack_12_field_type_1_sub_class_id : _GEN_5462; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5464 = _GEN_11433 & _GEN_10646 ? field_stack_12_field_type_2_sub_class_id : _GEN_5463; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5465 = _GEN_11433 & _GEN_10648 ? field_stack_12_field_type_3_sub_class_id : _GEN_5464; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5466 = _GEN_11433 & _GEN_10650 ? field_stack_12_field_type_4_sub_class_id : _GEN_5465; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5467 = _GEN_11433 & _GEN_10652 ? field_stack_12_field_type_5_sub_class_id : _GEN_5466; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5468 = _GEN_11433 & _GEN_10654 ? field_stack_12_field_type_6_sub_class_id : _GEN_5467; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5469 = _GEN_11433 & _GEN_10656 ? field_stack_12_field_type_7_sub_class_id : _GEN_5468; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5470 = _GEN_11433 & _GEN_10658 ? field_stack_12_field_type_8_sub_class_id : _GEN_5469; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5471 = _GEN_11433 & _GEN_10660 ? field_stack_12_field_type_9_sub_class_id : _GEN_5470; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5472 = _GEN_11433 & _GEN_10662 ? field_stack_12_field_type_10_sub_class_id : _GEN_5471; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5473 = _GEN_11433 & _GEN_10664 ? field_stack_12_field_type_11_sub_class_id : _GEN_5472; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5474 = _GEN_11433 & _GEN_10666 ? field_stack_12_field_type_12_sub_class_id : _GEN_5473; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5475 = _GEN_11433 & _GEN_10668 ? field_stack_12_field_type_13_sub_class_id : _GEN_5474; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5476 = _GEN_11433 & _GEN_10670 ? field_stack_12_field_type_14_sub_class_id : _GEN_5475; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5477 = _GEN_11433 & _GEN_10672 ? field_stack_12_field_type_15_sub_class_id : _GEN_5476; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5478 = _GEN_11433 & _GEN_10674 ? field_stack_12_field_type_16_sub_class_id : _GEN_5477; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5479 = _GEN_11433 & _GEN_10676 ? field_stack_12_field_type_17_sub_class_id : _GEN_5478; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5480 = _GEN_11433 & _GEN_10678 ? field_stack_12_field_type_18_sub_class_id : _GEN_5479; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5481 = _GEN_11433 & _GEN_10680 ? field_stack_12_field_type_19_sub_class_id : _GEN_5480; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5482 = _GEN_11433 & _GEN_10682 ? field_stack_12_field_type_20_sub_class_id : _GEN_5481; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5483 = _GEN_11433 & _GEN_10684 ? field_stack_12_field_type_21_sub_class_id : _GEN_5482; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5484 = _GEN_11433 & _GEN_10686 ? field_stack_12_field_type_22_sub_class_id : _GEN_5483; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5485 = _GEN_11433 & _GEN_10688 ? field_stack_12_field_type_23_sub_class_id : _GEN_5484; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5486 = _GEN_11433 & _GEN_10690 ? field_stack_12_field_type_24_sub_class_id : _GEN_5485; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5487 = _GEN_11433 & _GEN_10692 ? field_stack_12_field_type_25_sub_class_id : _GEN_5486; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5488 = _GEN_11433 & _GEN_10694 ? field_stack_12_field_type_26_sub_class_id : _GEN_5487; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5489 = _GEN_11433 & _GEN_10696 ? field_stack_12_field_type_27_sub_class_id : _GEN_5488; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5490 = _GEN_11433 & _GEN_10698 ? field_stack_12_field_type_28_sub_class_id : _GEN_5489; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5491 = _GEN_11433 & _GEN_10700 ? field_stack_12_field_type_29_sub_class_id : _GEN_5490; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5492 = _GEN_11433 & _GEN_10702 ? field_stack_12_field_type_30_sub_class_id : _GEN_5491; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5493 = _GEN_11433 & _GEN_10704 ? field_stack_12_field_type_31_sub_class_id : _GEN_5492; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5494 = _GEN_11433 & _GEN_10706 ? field_stack_12_field_type_32_sub_class_id : _GEN_5493; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5495 = _GEN_11499 & _GEN_10708 ? field_stack_13_field_type_0_sub_class_id : _GEN_5494; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5496 = _GEN_11499 & _GEN_10644 ? field_stack_13_field_type_1_sub_class_id : _GEN_5495; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5497 = _GEN_11499 & _GEN_10646 ? field_stack_13_field_type_2_sub_class_id : _GEN_5496; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5498 = _GEN_11499 & _GEN_10648 ? field_stack_13_field_type_3_sub_class_id : _GEN_5497; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5499 = _GEN_11499 & _GEN_10650 ? field_stack_13_field_type_4_sub_class_id : _GEN_5498; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5500 = _GEN_11499 & _GEN_10652 ? field_stack_13_field_type_5_sub_class_id : _GEN_5499; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5501 = _GEN_11499 & _GEN_10654 ? field_stack_13_field_type_6_sub_class_id : _GEN_5500; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5502 = _GEN_11499 & _GEN_10656 ? field_stack_13_field_type_7_sub_class_id : _GEN_5501; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5503 = _GEN_11499 & _GEN_10658 ? field_stack_13_field_type_8_sub_class_id : _GEN_5502; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5504 = _GEN_11499 & _GEN_10660 ? field_stack_13_field_type_9_sub_class_id : _GEN_5503; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5505 = _GEN_11499 & _GEN_10662 ? field_stack_13_field_type_10_sub_class_id : _GEN_5504; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5506 = _GEN_11499 & _GEN_10664 ? field_stack_13_field_type_11_sub_class_id : _GEN_5505; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5507 = _GEN_11499 & _GEN_10666 ? field_stack_13_field_type_12_sub_class_id : _GEN_5506; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5508 = _GEN_11499 & _GEN_10668 ? field_stack_13_field_type_13_sub_class_id : _GEN_5507; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5509 = _GEN_11499 & _GEN_10670 ? field_stack_13_field_type_14_sub_class_id : _GEN_5508; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5510 = _GEN_11499 & _GEN_10672 ? field_stack_13_field_type_15_sub_class_id : _GEN_5509; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5511 = _GEN_11499 & _GEN_10674 ? field_stack_13_field_type_16_sub_class_id : _GEN_5510; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5512 = _GEN_11499 & _GEN_10676 ? field_stack_13_field_type_17_sub_class_id : _GEN_5511; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5513 = _GEN_11499 & _GEN_10678 ? field_stack_13_field_type_18_sub_class_id : _GEN_5512; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5514 = _GEN_11499 & _GEN_10680 ? field_stack_13_field_type_19_sub_class_id : _GEN_5513; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5515 = _GEN_11499 & _GEN_10682 ? field_stack_13_field_type_20_sub_class_id : _GEN_5514; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5516 = _GEN_11499 & _GEN_10684 ? field_stack_13_field_type_21_sub_class_id : _GEN_5515; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5517 = _GEN_11499 & _GEN_10686 ? field_stack_13_field_type_22_sub_class_id : _GEN_5516; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5518 = _GEN_11499 & _GEN_10688 ? field_stack_13_field_type_23_sub_class_id : _GEN_5517; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5519 = _GEN_11499 & _GEN_10690 ? field_stack_13_field_type_24_sub_class_id : _GEN_5518; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5520 = _GEN_11499 & _GEN_10692 ? field_stack_13_field_type_25_sub_class_id : _GEN_5519; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5521 = _GEN_11499 & _GEN_10694 ? field_stack_13_field_type_26_sub_class_id : _GEN_5520; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5522 = _GEN_11499 & _GEN_10696 ? field_stack_13_field_type_27_sub_class_id : _GEN_5521; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5523 = _GEN_11499 & _GEN_10698 ? field_stack_13_field_type_28_sub_class_id : _GEN_5522; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5524 = _GEN_11499 & _GEN_10700 ? field_stack_13_field_type_29_sub_class_id : _GEN_5523; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5525 = _GEN_11499 & _GEN_10702 ? field_stack_13_field_type_30_sub_class_id : _GEN_5524; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5526 = _GEN_11499 & _GEN_10704 ? field_stack_13_field_type_31_sub_class_id : _GEN_5525; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5527 = _GEN_11499 & _GEN_10706 ? field_stack_13_field_type_32_sub_class_id : _GEN_5526; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5528 = _GEN_11565 & _GEN_10708 ? field_stack_14_field_type_0_sub_class_id : _GEN_5527; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5529 = _GEN_11565 & _GEN_10644 ? field_stack_14_field_type_1_sub_class_id : _GEN_5528; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5530 = _GEN_11565 & _GEN_10646 ? field_stack_14_field_type_2_sub_class_id : _GEN_5529; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5531 = _GEN_11565 & _GEN_10648 ? field_stack_14_field_type_3_sub_class_id : _GEN_5530; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5532 = _GEN_11565 & _GEN_10650 ? field_stack_14_field_type_4_sub_class_id : _GEN_5531; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5533 = _GEN_11565 & _GEN_10652 ? field_stack_14_field_type_5_sub_class_id : _GEN_5532; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5534 = _GEN_11565 & _GEN_10654 ? field_stack_14_field_type_6_sub_class_id : _GEN_5533; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5535 = _GEN_11565 & _GEN_10656 ? field_stack_14_field_type_7_sub_class_id : _GEN_5534; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5536 = _GEN_11565 & _GEN_10658 ? field_stack_14_field_type_8_sub_class_id : _GEN_5535; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5537 = _GEN_11565 & _GEN_10660 ? field_stack_14_field_type_9_sub_class_id : _GEN_5536; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5538 = _GEN_11565 & _GEN_10662 ? field_stack_14_field_type_10_sub_class_id : _GEN_5537; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5539 = _GEN_11565 & _GEN_10664 ? field_stack_14_field_type_11_sub_class_id : _GEN_5538; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5540 = _GEN_11565 & _GEN_10666 ? field_stack_14_field_type_12_sub_class_id : _GEN_5539; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5541 = _GEN_11565 & _GEN_10668 ? field_stack_14_field_type_13_sub_class_id : _GEN_5540; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5542 = _GEN_11565 & _GEN_10670 ? field_stack_14_field_type_14_sub_class_id : _GEN_5541; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5543 = _GEN_11565 & _GEN_10672 ? field_stack_14_field_type_15_sub_class_id : _GEN_5542; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5544 = _GEN_11565 & _GEN_10674 ? field_stack_14_field_type_16_sub_class_id : _GEN_5543; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5545 = _GEN_11565 & _GEN_10676 ? field_stack_14_field_type_17_sub_class_id : _GEN_5544; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5546 = _GEN_11565 & _GEN_10678 ? field_stack_14_field_type_18_sub_class_id : _GEN_5545; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5547 = _GEN_11565 & _GEN_10680 ? field_stack_14_field_type_19_sub_class_id : _GEN_5546; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5548 = _GEN_11565 & _GEN_10682 ? field_stack_14_field_type_20_sub_class_id : _GEN_5547; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5549 = _GEN_11565 & _GEN_10684 ? field_stack_14_field_type_21_sub_class_id : _GEN_5548; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5550 = _GEN_11565 & _GEN_10686 ? field_stack_14_field_type_22_sub_class_id : _GEN_5549; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5551 = _GEN_11565 & _GEN_10688 ? field_stack_14_field_type_23_sub_class_id : _GEN_5550; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5552 = _GEN_11565 & _GEN_10690 ? field_stack_14_field_type_24_sub_class_id : _GEN_5551; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5553 = _GEN_11565 & _GEN_10692 ? field_stack_14_field_type_25_sub_class_id : _GEN_5552; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5554 = _GEN_11565 & _GEN_10694 ? field_stack_14_field_type_26_sub_class_id : _GEN_5553; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5555 = _GEN_11565 & _GEN_10696 ? field_stack_14_field_type_27_sub_class_id : _GEN_5554; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5556 = _GEN_11565 & _GEN_10698 ? field_stack_14_field_type_28_sub_class_id : _GEN_5555; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5557 = _GEN_11565 & _GEN_10700 ? field_stack_14_field_type_29_sub_class_id : _GEN_5556; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5558 = _GEN_11565 & _GEN_10702 ? field_stack_14_field_type_30_sub_class_id : _GEN_5557; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5559 = _GEN_11565 & _GEN_10704 ? field_stack_14_field_type_31_sub_class_id : _GEN_5558; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [15:0] _GEN_5560 = _GEN_11565 & _GEN_10706 ? field_stack_14_field_type_32_sub_class_id : _GEN_5559; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5562 = _GEN_10643 & _GEN_10644 ? field_stack_0_field_type_1_is_repeated :
    field_stack_0_field_type_0_is_repeated; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5563 = _GEN_10643 & _GEN_10646 ? field_stack_0_field_type_2_is_repeated : _GEN_5562; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5564 = _GEN_10643 & _GEN_10648 ? field_stack_0_field_type_3_is_repeated : _GEN_5563; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5565 = _GEN_10643 & _GEN_10650 ? field_stack_0_field_type_4_is_repeated : _GEN_5564; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5566 = _GEN_10643 & _GEN_10652 ? field_stack_0_field_type_5_is_repeated : _GEN_5565; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5567 = _GEN_10643 & _GEN_10654 ? field_stack_0_field_type_6_is_repeated : _GEN_5566; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5568 = _GEN_10643 & _GEN_10656 ? field_stack_0_field_type_7_is_repeated : _GEN_5567; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5569 = _GEN_10643 & _GEN_10658 ? field_stack_0_field_type_8_is_repeated : _GEN_5568; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5570 = _GEN_10643 & _GEN_10660 ? field_stack_0_field_type_9_is_repeated : _GEN_5569; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5571 = _GEN_10643 & _GEN_10662 ? field_stack_0_field_type_10_is_repeated : _GEN_5570; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5572 = _GEN_10643 & _GEN_10664 ? field_stack_0_field_type_11_is_repeated : _GEN_5571; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5573 = _GEN_10643 & _GEN_10666 ? field_stack_0_field_type_12_is_repeated : _GEN_5572; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5574 = _GEN_10643 & _GEN_10668 ? field_stack_0_field_type_13_is_repeated : _GEN_5573; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5575 = _GEN_10643 & _GEN_10670 ? field_stack_0_field_type_14_is_repeated : _GEN_5574; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5576 = _GEN_10643 & _GEN_10672 ? field_stack_0_field_type_15_is_repeated : _GEN_5575; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5577 = _GEN_10643 & _GEN_10674 ? field_stack_0_field_type_16_is_repeated : _GEN_5576; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5578 = _GEN_10643 & _GEN_10676 ? field_stack_0_field_type_17_is_repeated : _GEN_5577; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5579 = _GEN_10643 & _GEN_10678 ? field_stack_0_field_type_18_is_repeated : _GEN_5578; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5580 = _GEN_10643 & _GEN_10680 ? field_stack_0_field_type_19_is_repeated : _GEN_5579; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5581 = _GEN_10643 & _GEN_10682 ? field_stack_0_field_type_20_is_repeated : _GEN_5580; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5582 = _GEN_10643 & _GEN_10684 ? field_stack_0_field_type_21_is_repeated : _GEN_5581; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5583 = _GEN_10643 & _GEN_10686 ? field_stack_0_field_type_22_is_repeated : _GEN_5582; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5584 = _GEN_10643 & _GEN_10688 ? field_stack_0_field_type_23_is_repeated : _GEN_5583; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5585 = _GEN_10643 & _GEN_10690 ? field_stack_0_field_type_24_is_repeated : _GEN_5584; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5586 = _GEN_10643 & _GEN_10692 ? field_stack_0_field_type_25_is_repeated : _GEN_5585; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5587 = _GEN_10643 & _GEN_10694 ? field_stack_0_field_type_26_is_repeated : _GEN_5586; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5588 = _GEN_10643 & _GEN_10696 ? field_stack_0_field_type_27_is_repeated : _GEN_5587; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5589 = _GEN_10643 & _GEN_10698 ? field_stack_0_field_type_28_is_repeated : _GEN_5588; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5590 = _GEN_10643 & _GEN_10700 ? field_stack_0_field_type_29_is_repeated : _GEN_5589; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5591 = _GEN_10643 & _GEN_10702 ? field_stack_0_field_type_30_is_repeated : _GEN_5590; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5592 = _GEN_10643 & _GEN_10704 ? field_stack_0_field_type_31_is_repeated : _GEN_5591; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5593 = _GEN_10643 & _GEN_10706 ? field_stack_0_field_type_32_is_repeated : _GEN_5592; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5594 = _GEN_10707 & _GEN_10708 ? field_stack_1_field_type_0_is_repeated : _GEN_5593; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5595 = _GEN_10707 & _GEN_10644 ? field_stack_1_field_type_1_is_repeated : _GEN_5594; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5596 = _GEN_10707 & _GEN_10646 ? field_stack_1_field_type_2_is_repeated : _GEN_5595; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5597 = _GEN_10707 & _GEN_10648 ? field_stack_1_field_type_3_is_repeated : _GEN_5596; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5598 = _GEN_10707 & _GEN_10650 ? field_stack_1_field_type_4_is_repeated : _GEN_5597; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5599 = _GEN_10707 & _GEN_10652 ? field_stack_1_field_type_5_is_repeated : _GEN_5598; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5600 = _GEN_10707 & _GEN_10654 ? field_stack_1_field_type_6_is_repeated : _GEN_5599; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5601 = _GEN_10707 & _GEN_10656 ? field_stack_1_field_type_7_is_repeated : _GEN_5600; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5602 = _GEN_10707 & _GEN_10658 ? field_stack_1_field_type_8_is_repeated : _GEN_5601; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5603 = _GEN_10707 & _GEN_10660 ? field_stack_1_field_type_9_is_repeated : _GEN_5602; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5604 = _GEN_10707 & _GEN_10662 ? field_stack_1_field_type_10_is_repeated : _GEN_5603; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5605 = _GEN_10707 & _GEN_10664 ? field_stack_1_field_type_11_is_repeated : _GEN_5604; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5606 = _GEN_10707 & _GEN_10666 ? field_stack_1_field_type_12_is_repeated : _GEN_5605; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5607 = _GEN_10707 & _GEN_10668 ? field_stack_1_field_type_13_is_repeated : _GEN_5606; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5608 = _GEN_10707 & _GEN_10670 ? field_stack_1_field_type_14_is_repeated : _GEN_5607; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5609 = _GEN_10707 & _GEN_10672 ? field_stack_1_field_type_15_is_repeated : _GEN_5608; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5610 = _GEN_10707 & _GEN_10674 ? field_stack_1_field_type_16_is_repeated : _GEN_5609; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5611 = _GEN_10707 & _GEN_10676 ? field_stack_1_field_type_17_is_repeated : _GEN_5610; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5612 = _GEN_10707 & _GEN_10678 ? field_stack_1_field_type_18_is_repeated : _GEN_5611; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5613 = _GEN_10707 & _GEN_10680 ? field_stack_1_field_type_19_is_repeated : _GEN_5612; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5614 = _GEN_10707 & _GEN_10682 ? field_stack_1_field_type_20_is_repeated : _GEN_5613; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5615 = _GEN_10707 & _GEN_10684 ? field_stack_1_field_type_21_is_repeated : _GEN_5614; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5616 = _GEN_10707 & _GEN_10686 ? field_stack_1_field_type_22_is_repeated : _GEN_5615; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5617 = _GEN_10707 & _GEN_10688 ? field_stack_1_field_type_23_is_repeated : _GEN_5616; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5618 = _GEN_10707 & _GEN_10690 ? field_stack_1_field_type_24_is_repeated : _GEN_5617; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5619 = _GEN_10707 & _GEN_10692 ? field_stack_1_field_type_25_is_repeated : _GEN_5618; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5620 = _GEN_10707 & _GEN_10694 ? field_stack_1_field_type_26_is_repeated : _GEN_5619; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5621 = _GEN_10707 & _GEN_10696 ? field_stack_1_field_type_27_is_repeated : _GEN_5620; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5622 = _GEN_10707 & _GEN_10698 ? field_stack_1_field_type_28_is_repeated : _GEN_5621; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5623 = _GEN_10707 & _GEN_10700 ? field_stack_1_field_type_29_is_repeated : _GEN_5622; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5624 = _GEN_10707 & _GEN_10702 ? field_stack_1_field_type_30_is_repeated : _GEN_5623; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5625 = _GEN_10707 & _GEN_10704 ? field_stack_1_field_type_31_is_repeated : _GEN_5624; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5626 = _GEN_10707 & _GEN_10706 ? field_stack_1_field_type_32_is_repeated : _GEN_5625; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5627 = _GEN_10773 & _GEN_10708 ? field_stack_2_field_type_0_is_repeated : _GEN_5626; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5628 = _GEN_10773 & _GEN_10644 ? field_stack_2_field_type_1_is_repeated : _GEN_5627; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5629 = _GEN_10773 & _GEN_10646 ? field_stack_2_field_type_2_is_repeated : _GEN_5628; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5630 = _GEN_10773 & _GEN_10648 ? field_stack_2_field_type_3_is_repeated : _GEN_5629; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5631 = _GEN_10773 & _GEN_10650 ? field_stack_2_field_type_4_is_repeated : _GEN_5630; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5632 = _GEN_10773 & _GEN_10652 ? field_stack_2_field_type_5_is_repeated : _GEN_5631; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5633 = _GEN_10773 & _GEN_10654 ? field_stack_2_field_type_6_is_repeated : _GEN_5632; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5634 = _GEN_10773 & _GEN_10656 ? field_stack_2_field_type_7_is_repeated : _GEN_5633; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5635 = _GEN_10773 & _GEN_10658 ? field_stack_2_field_type_8_is_repeated : _GEN_5634; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5636 = _GEN_10773 & _GEN_10660 ? field_stack_2_field_type_9_is_repeated : _GEN_5635; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5637 = _GEN_10773 & _GEN_10662 ? field_stack_2_field_type_10_is_repeated : _GEN_5636; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5638 = _GEN_10773 & _GEN_10664 ? field_stack_2_field_type_11_is_repeated : _GEN_5637; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5639 = _GEN_10773 & _GEN_10666 ? field_stack_2_field_type_12_is_repeated : _GEN_5638; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5640 = _GEN_10773 & _GEN_10668 ? field_stack_2_field_type_13_is_repeated : _GEN_5639; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5641 = _GEN_10773 & _GEN_10670 ? field_stack_2_field_type_14_is_repeated : _GEN_5640; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5642 = _GEN_10773 & _GEN_10672 ? field_stack_2_field_type_15_is_repeated : _GEN_5641; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5643 = _GEN_10773 & _GEN_10674 ? field_stack_2_field_type_16_is_repeated : _GEN_5642; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5644 = _GEN_10773 & _GEN_10676 ? field_stack_2_field_type_17_is_repeated : _GEN_5643; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5645 = _GEN_10773 & _GEN_10678 ? field_stack_2_field_type_18_is_repeated : _GEN_5644; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5646 = _GEN_10773 & _GEN_10680 ? field_stack_2_field_type_19_is_repeated : _GEN_5645; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5647 = _GEN_10773 & _GEN_10682 ? field_stack_2_field_type_20_is_repeated : _GEN_5646; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5648 = _GEN_10773 & _GEN_10684 ? field_stack_2_field_type_21_is_repeated : _GEN_5647; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5649 = _GEN_10773 & _GEN_10686 ? field_stack_2_field_type_22_is_repeated : _GEN_5648; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5650 = _GEN_10773 & _GEN_10688 ? field_stack_2_field_type_23_is_repeated : _GEN_5649; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5651 = _GEN_10773 & _GEN_10690 ? field_stack_2_field_type_24_is_repeated : _GEN_5650; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5652 = _GEN_10773 & _GEN_10692 ? field_stack_2_field_type_25_is_repeated : _GEN_5651; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5653 = _GEN_10773 & _GEN_10694 ? field_stack_2_field_type_26_is_repeated : _GEN_5652; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5654 = _GEN_10773 & _GEN_10696 ? field_stack_2_field_type_27_is_repeated : _GEN_5653; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5655 = _GEN_10773 & _GEN_10698 ? field_stack_2_field_type_28_is_repeated : _GEN_5654; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5656 = _GEN_10773 & _GEN_10700 ? field_stack_2_field_type_29_is_repeated : _GEN_5655; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5657 = _GEN_10773 & _GEN_10702 ? field_stack_2_field_type_30_is_repeated : _GEN_5656; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5658 = _GEN_10773 & _GEN_10704 ? field_stack_2_field_type_31_is_repeated : _GEN_5657; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5659 = _GEN_10773 & _GEN_10706 ? field_stack_2_field_type_32_is_repeated : _GEN_5658; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5660 = _GEN_10839 & _GEN_10708 ? field_stack_3_field_type_0_is_repeated : _GEN_5659; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5661 = _GEN_10839 & _GEN_10644 ? field_stack_3_field_type_1_is_repeated : _GEN_5660; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5662 = _GEN_10839 & _GEN_10646 ? field_stack_3_field_type_2_is_repeated : _GEN_5661; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5663 = _GEN_10839 & _GEN_10648 ? field_stack_3_field_type_3_is_repeated : _GEN_5662; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5664 = _GEN_10839 & _GEN_10650 ? field_stack_3_field_type_4_is_repeated : _GEN_5663; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5665 = _GEN_10839 & _GEN_10652 ? field_stack_3_field_type_5_is_repeated : _GEN_5664; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5666 = _GEN_10839 & _GEN_10654 ? field_stack_3_field_type_6_is_repeated : _GEN_5665; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5667 = _GEN_10839 & _GEN_10656 ? field_stack_3_field_type_7_is_repeated : _GEN_5666; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5668 = _GEN_10839 & _GEN_10658 ? field_stack_3_field_type_8_is_repeated : _GEN_5667; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5669 = _GEN_10839 & _GEN_10660 ? field_stack_3_field_type_9_is_repeated : _GEN_5668; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5670 = _GEN_10839 & _GEN_10662 ? field_stack_3_field_type_10_is_repeated : _GEN_5669; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5671 = _GEN_10839 & _GEN_10664 ? field_stack_3_field_type_11_is_repeated : _GEN_5670; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5672 = _GEN_10839 & _GEN_10666 ? field_stack_3_field_type_12_is_repeated : _GEN_5671; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5673 = _GEN_10839 & _GEN_10668 ? field_stack_3_field_type_13_is_repeated : _GEN_5672; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5674 = _GEN_10839 & _GEN_10670 ? field_stack_3_field_type_14_is_repeated : _GEN_5673; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5675 = _GEN_10839 & _GEN_10672 ? field_stack_3_field_type_15_is_repeated : _GEN_5674; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5676 = _GEN_10839 & _GEN_10674 ? field_stack_3_field_type_16_is_repeated : _GEN_5675; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5677 = _GEN_10839 & _GEN_10676 ? field_stack_3_field_type_17_is_repeated : _GEN_5676; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5678 = _GEN_10839 & _GEN_10678 ? field_stack_3_field_type_18_is_repeated : _GEN_5677; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5679 = _GEN_10839 & _GEN_10680 ? field_stack_3_field_type_19_is_repeated : _GEN_5678; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5680 = _GEN_10839 & _GEN_10682 ? field_stack_3_field_type_20_is_repeated : _GEN_5679; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5681 = _GEN_10839 & _GEN_10684 ? field_stack_3_field_type_21_is_repeated : _GEN_5680; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5682 = _GEN_10839 & _GEN_10686 ? field_stack_3_field_type_22_is_repeated : _GEN_5681; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5683 = _GEN_10839 & _GEN_10688 ? field_stack_3_field_type_23_is_repeated : _GEN_5682; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5684 = _GEN_10839 & _GEN_10690 ? field_stack_3_field_type_24_is_repeated : _GEN_5683; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5685 = _GEN_10839 & _GEN_10692 ? field_stack_3_field_type_25_is_repeated : _GEN_5684; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5686 = _GEN_10839 & _GEN_10694 ? field_stack_3_field_type_26_is_repeated : _GEN_5685; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5687 = _GEN_10839 & _GEN_10696 ? field_stack_3_field_type_27_is_repeated : _GEN_5686; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5688 = _GEN_10839 & _GEN_10698 ? field_stack_3_field_type_28_is_repeated : _GEN_5687; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5689 = _GEN_10839 & _GEN_10700 ? field_stack_3_field_type_29_is_repeated : _GEN_5688; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5690 = _GEN_10839 & _GEN_10702 ? field_stack_3_field_type_30_is_repeated : _GEN_5689; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5691 = _GEN_10839 & _GEN_10704 ? field_stack_3_field_type_31_is_repeated : _GEN_5690; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5692 = _GEN_10839 & _GEN_10706 ? field_stack_3_field_type_32_is_repeated : _GEN_5691; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5693 = _GEN_10905 & _GEN_10708 ? field_stack_4_field_type_0_is_repeated : _GEN_5692; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5694 = _GEN_10905 & _GEN_10644 ? field_stack_4_field_type_1_is_repeated : _GEN_5693; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5695 = _GEN_10905 & _GEN_10646 ? field_stack_4_field_type_2_is_repeated : _GEN_5694; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5696 = _GEN_10905 & _GEN_10648 ? field_stack_4_field_type_3_is_repeated : _GEN_5695; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5697 = _GEN_10905 & _GEN_10650 ? field_stack_4_field_type_4_is_repeated : _GEN_5696; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5698 = _GEN_10905 & _GEN_10652 ? field_stack_4_field_type_5_is_repeated : _GEN_5697; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5699 = _GEN_10905 & _GEN_10654 ? field_stack_4_field_type_6_is_repeated : _GEN_5698; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5700 = _GEN_10905 & _GEN_10656 ? field_stack_4_field_type_7_is_repeated : _GEN_5699; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5701 = _GEN_10905 & _GEN_10658 ? field_stack_4_field_type_8_is_repeated : _GEN_5700; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5702 = _GEN_10905 & _GEN_10660 ? field_stack_4_field_type_9_is_repeated : _GEN_5701; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5703 = _GEN_10905 & _GEN_10662 ? field_stack_4_field_type_10_is_repeated : _GEN_5702; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5704 = _GEN_10905 & _GEN_10664 ? field_stack_4_field_type_11_is_repeated : _GEN_5703; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5705 = _GEN_10905 & _GEN_10666 ? field_stack_4_field_type_12_is_repeated : _GEN_5704; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5706 = _GEN_10905 & _GEN_10668 ? field_stack_4_field_type_13_is_repeated : _GEN_5705; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5707 = _GEN_10905 & _GEN_10670 ? field_stack_4_field_type_14_is_repeated : _GEN_5706; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5708 = _GEN_10905 & _GEN_10672 ? field_stack_4_field_type_15_is_repeated : _GEN_5707; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5709 = _GEN_10905 & _GEN_10674 ? field_stack_4_field_type_16_is_repeated : _GEN_5708; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5710 = _GEN_10905 & _GEN_10676 ? field_stack_4_field_type_17_is_repeated : _GEN_5709; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5711 = _GEN_10905 & _GEN_10678 ? field_stack_4_field_type_18_is_repeated : _GEN_5710; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5712 = _GEN_10905 & _GEN_10680 ? field_stack_4_field_type_19_is_repeated : _GEN_5711; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5713 = _GEN_10905 & _GEN_10682 ? field_stack_4_field_type_20_is_repeated : _GEN_5712; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5714 = _GEN_10905 & _GEN_10684 ? field_stack_4_field_type_21_is_repeated : _GEN_5713; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5715 = _GEN_10905 & _GEN_10686 ? field_stack_4_field_type_22_is_repeated : _GEN_5714; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5716 = _GEN_10905 & _GEN_10688 ? field_stack_4_field_type_23_is_repeated : _GEN_5715; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5717 = _GEN_10905 & _GEN_10690 ? field_stack_4_field_type_24_is_repeated : _GEN_5716; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5718 = _GEN_10905 & _GEN_10692 ? field_stack_4_field_type_25_is_repeated : _GEN_5717; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5719 = _GEN_10905 & _GEN_10694 ? field_stack_4_field_type_26_is_repeated : _GEN_5718; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5720 = _GEN_10905 & _GEN_10696 ? field_stack_4_field_type_27_is_repeated : _GEN_5719; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5721 = _GEN_10905 & _GEN_10698 ? field_stack_4_field_type_28_is_repeated : _GEN_5720; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5722 = _GEN_10905 & _GEN_10700 ? field_stack_4_field_type_29_is_repeated : _GEN_5721; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5723 = _GEN_10905 & _GEN_10702 ? field_stack_4_field_type_30_is_repeated : _GEN_5722; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5724 = _GEN_10905 & _GEN_10704 ? field_stack_4_field_type_31_is_repeated : _GEN_5723; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5725 = _GEN_10905 & _GEN_10706 ? field_stack_4_field_type_32_is_repeated : _GEN_5724; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5726 = _GEN_10971 & _GEN_10708 ? field_stack_5_field_type_0_is_repeated : _GEN_5725; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5727 = _GEN_10971 & _GEN_10644 ? field_stack_5_field_type_1_is_repeated : _GEN_5726; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5728 = _GEN_10971 & _GEN_10646 ? field_stack_5_field_type_2_is_repeated : _GEN_5727; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5729 = _GEN_10971 & _GEN_10648 ? field_stack_5_field_type_3_is_repeated : _GEN_5728; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5730 = _GEN_10971 & _GEN_10650 ? field_stack_5_field_type_4_is_repeated : _GEN_5729; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5731 = _GEN_10971 & _GEN_10652 ? field_stack_5_field_type_5_is_repeated : _GEN_5730; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5732 = _GEN_10971 & _GEN_10654 ? field_stack_5_field_type_6_is_repeated : _GEN_5731; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5733 = _GEN_10971 & _GEN_10656 ? field_stack_5_field_type_7_is_repeated : _GEN_5732; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5734 = _GEN_10971 & _GEN_10658 ? field_stack_5_field_type_8_is_repeated : _GEN_5733; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5735 = _GEN_10971 & _GEN_10660 ? field_stack_5_field_type_9_is_repeated : _GEN_5734; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5736 = _GEN_10971 & _GEN_10662 ? field_stack_5_field_type_10_is_repeated : _GEN_5735; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5737 = _GEN_10971 & _GEN_10664 ? field_stack_5_field_type_11_is_repeated : _GEN_5736; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5738 = _GEN_10971 & _GEN_10666 ? field_stack_5_field_type_12_is_repeated : _GEN_5737; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5739 = _GEN_10971 & _GEN_10668 ? field_stack_5_field_type_13_is_repeated : _GEN_5738; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5740 = _GEN_10971 & _GEN_10670 ? field_stack_5_field_type_14_is_repeated : _GEN_5739; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5741 = _GEN_10971 & _GEN_10672 ? field_stack_5_field_type_15_is_repeated : _GEN_5740; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5742 = _GEN_10971 & _GEN_10674 ? field_stack_5_field_type_16_is_repeated : _GEN_5741; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5743 = _GEN_10971 & _GEN_10676 ? field_stack_5_field_type_17_is_repeated : _GEN_5742; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5744 = _GEN_10971 & _GEN_10678 ? field_stack_5_field_type_18_is_repeated : _GEN_5743; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5745 = _GEN_10971 & _GEN_10680 ? field_stack_5_field_type_19_is_repeated : _GEN_5744; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5746 = _GEN_10971 & _GEN_10682 ? field_stack_5_field_type_20_is_repeated : _GEN_5745; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5747 = _GEN_10971 & _GEN_10684 ? field_stack_5_field_type_21_is_repeated : _GEN_5746; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5748 = _GEN_10971 & _GEN_10686 ? field_stack_5_field_type_22_is_repeated : _GEN_5747; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5749 = _GEN_10971 & _GEN_10688 ? field_stack_5_field_type_23_is_repeated : _GEN_5748; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5750 = _GEN_10971 & _GEN_10690 ? field_stack_5_field_type_24_is_repeated : _GEN_5749; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5751 = _GEN_10971 & _GEN_10692 ? field_stack_5_field_type_25_is_repeated : _GEN_5750; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5752 = _GEN_10971 & _GEN_10694 ? field_stack_5_field_type_26_is_repeated : _GEN_5751; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5753 = _GEN_10971 & _GEN_10696 ? field_stack_5_field_type_27_is_repeated : _GEN_5752; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5754 = _GEN_10971 & _GEN_10698 ? field_stack_5_field_type_28_is_repeated : _GEN_5753; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5755 = _GEN_10971 & _GEN_10700 ? field_stack_5_field_type_29_is_repeated : _GEN_5754; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5756 = _GEN_10971 & _GEN_10702 ? field_stack_5_field_type_30_is_repeated : _GEN_5755; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5757 = _GEN_10971 & _GEN_10704 ? field_stack_5_field_type_31_is_repeated : _GEN_5756; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5758 = _GEN_10971 & _GEN_10706 ? field_stack_5_field_type_32_is_repeated : _GEN_5757; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5759 = _GEN_11037 & _GEN_10708 ? field_stack_6_field_type_0_is_repeated : _GEN_5758; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5760 = _GEN_11037 & _GEN_10644 ? field_stack_6_field_type_1_is_repeated : _GEN_5759; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5761 = _GEN_11037 & _GEN_10646 ? field_stack_6_field_type_2_is_repeated : _GEN_5760; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5762 = _GEN_11037 & _GEN_10648 ? field_stack_6_field_type_3_is_repeated : _GEN_5761; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5763 = _GEN_11037 & _GEN_10650 ? field_stack_6_field_type_4_is_repeated : _GEN_5762; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5764 = _GEN_11037 & _GEN_10652 ? field_stack_6_field_type_5_is_repeated : _GEN_5763; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5765 = _GEN_11037 & _GEN_10654 ? field_stack_6_field_type_6_is_repeated : _GEN_5764; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5766 = _GEN_11037 & _GEN_10656 ? field_stack_6_field_type_7_is_repeated : _GEN_5765; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5767 = _GEN_11037 & _GEN_10658 ? field_stack_6_field_type_8_is_repeated : _GEN_5766; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5768 = _GEN_11037 & _GEN_10660 ? field_stack_6_field_type_9_is_repeated : _GEN_5767; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5769 = _GEN_11037 & _GEN_10662 ? field_stack_6_field_type_10_is_repeated : _GEN_5768; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5770 = _GEN_11037 & _GEN_10664 ? field_stack_6_field_type_11_is_repeated : _GEN_5769; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5771 = _GEN_11037 & _GEN_10666 ? field_stack_6_field_type_12_is_repeated : _GEN_5770; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5772 = _GEN_11037 & _GEN_10668 ? field_stack_6_field_type_13_is_repeated : _GEN_5771; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5773 = _GEN_11037 & _GEN_10670 ? field_stack_6_field_type_14_is_repeated : _GEN_5772; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5774 = _GEN_11037 & _GEN_10672 ? field_stack_6_field_type_15_is_repeated : _GEN_5773; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5775 = _GEN_11037 & _GEN_10674 ? field_stack_6_field_type_16_is_repeated : _GEN_5774; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5776 = _GEN_11037 & _GEN_10676 ? field_stack_6_field_type_17_is_repeated : _GEN_5775; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5777 = _GEN_11037 & _GEN_10678 ? field_stack_6_field_type_18_is_repeated : _GEN_5776; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5778 = _GEN_11037 & _GEN_10680 ? field_stack_6_field_type_19_is_repeated : _GEN_5777; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5779 = _GEN_11037 & _GEN_10682 ? field_stack_6_field_type_20_is_repeated : _GEN_5778; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5780 = _GEN_11037 & _GEN_10684 ? field_stack_6_field_type_21_is_repeated : _GEN_5779; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5781 = _GEN_11037 & _GEN_10686 ? field_stack_6_field_type_22_is_repeated : _GEN_5780; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5782 = _GEN_11037 & _GEN_10688 ? field_stack_6_field_type_23_is_repeated : _GEN_5781; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5783 = _GEN_11037 & _GEN_10690 ? field_stack_6_field_type_24_is_repeated : _GEN_5782; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5784 = _GEN_11037 & _GEN_10692 ? field_stack_6_field_type_25_is_repeated : _GEN_5783; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5785 = _GEN_11037 & _GEN_10694 ? field_stack_6_field_type_26_is_repeated : _GEN_5784; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5786 = _GEN_11037 & _GEN_10696 ? field_stack_6_field_type_27_is_repeated : _GEN_5785; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5787 = _GEN_11037 & _GEN_10698 ? field_stack_6_field_type_28_is_repeated : _GEN_5786; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5788 = _GEN_11037 & _GEN_10700 ? field_stack_6_field_type_29_is_repeated : _GEN_5787; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5789 = _GEN_11037 & _GEN_10702 ? field_stack_6_field_type_30_is_repeated : _GEN_5788; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5790 = _GEN_11037 & _GEN_10704 ? field_stack_6_field_type_31_is_repeated : _GEN_5789; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5791 = _GEN_11037 & _GEN_10706 ? field_stack_6_field_type_32_is_repeated : _GEN_5790; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5792 = _GEN_11103 & _GEN_10708 ? field_stack_7_field_type_0_is_repeated : _GEN_5791; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5793 = _GEN_11103 & _GEN_10644 ? field_stack_7_field_type_1_is_repeated : _GEN_5792; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5794 = _GEN_11103 & _GEN_10646 ? field_stack_7_field_type_2_is_repeated : _GEN_5793; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5795 = _GEN_11103 & _GEN_10648 ? field_stack_7_field_type_3_is_repeated : _GEN_5794; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5796 = _GEN_11103 & _GEN_10650 ? field_stack_7_field_type_4_is_repeated : _GEN_5795; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5797 = _GEN_11103 & _GEN_10652 ? field_stack_7_field_type_5_is_repeated : _GEN_5796; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5798 = _GEN_11103 & _GEN_10654 ? field_stack_7_field_type_6_is_repeated : _GEN_5797; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5799 = _GEN_11103 & _GEN_10656 ? field_stack_7_field_type_7_is_repeated : _GEN_5798; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5800 = _GEN_11103 & _GEN_10658 ? field_stack_7_field_type_8_is_repeated : _GEN_5799; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5801 = _GEN_11103 & _GEN_10660 ? field_stack_7_field_type_9_is_repeated : _GEN_5800; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5802 = _GEN_11103 & _GEN_10662 ? field_stack_7_field_type_10_is_repeated : _GEN_5801; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5803 = _GEN_11103 & _GEN_10664 ? field_stack_7_field_type_11_is_repeated : _GEN_5802; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5804 = _GEN_11103 & _GEN_10666 ? field_stack_7_field_type_12_is_repeated : _GEN_5803; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5805 = _GEN_11103 & _GEN_10668 ? field_stack_7_field_type_13_is_repeated : _GEN_5804; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5806 = _GEN_11103 & _GEN_10670 ? field_stack_7_field_type_14_is_repeated : _GEN_5805; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5807 = _GEN_11103 & _GEN_10672 ? field_stack_7_field_type_15_is_repeated : _GEN_5806; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5808 = _GEN_11103 & _GEN_10674 ? field_stack_7_field_type_16_is_repeated : _GEN_5807; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5809 = _GEN_11103 & _GEN_10676 ? field_stack_7_field_type_17_is_repeated : _GEN_5808; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5810 = _GEN_11103 & _GEN_10678 ? field_stack_7_field_type_18_is_repeated : _GEN_5809; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5811 = _GEN_11103 & _GEN_10680 ? field_stack_7_field_type_19_is_repeated : _GEN_5810; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5812 = _GEN_11103 & _GEN_10682 ? field_stack_7_field_type_20_is_repeated : _GEN_5811; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5813 = _GEN_11103 & _GEN_10684 ? field_stack_7_field_type_21_is_repeated : _GEN_5812; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5814 = _GEN_11103 & _GEN_10686 ? field_stack_7_field_type_22_is_repeated : _GEN_5813; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5815 = _GEN_11103 & _GEN_10688 ? field_stack_7_field_type_23_is_repeated : _GEN_5814; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5816 = _GEN_11103 & _GEN_10690 ? field_stack_7_field_type_24_is_repeated : _GEN_5815; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5817 = _GEN_11103 & _GEN_10692 ? field_stack_7_field_type_25_is_repeated : _GEN_5816; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5818 = _GEN_11103 & _GEN_10694 ? field_stack_7_field_type_26_is_repeated : _GEN_5817; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5819 = _GEN_11103 & _GEN_10696 ? field_stack_7_field_type_27_is_repeated : _GEN_5818; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5820 = _GEN_11103 & _GEN_10698 ? field_stack_7_field_type_28_is_repeated : _GEN_5819; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5821 = _GEN_11103 & _GEN_10700 ? field_stack_7_field_type_29_is_repeated : _GEN_5820; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5822 = _GEN_11103 & _GEN_10702 ? field_stack_7_field_type_30_is_repeated : _GEN_5821; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5823 = _GEN_11103 & _GEN_10704 ? field_stack_7_field_type_31_is_repeated : _GEN_5822; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5824 = _GEN_11103 & _GEN_10706 ? field_stack_7_field_type_32_is_repeated : _GEN_5823; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5825 = _GEN_11169 & _GEN_10708 ? field_stack_8_field_type_0_is_repeated : _GEN_5824; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5826 = _GEN_11169 & _GEN_10644 ? field_stack_8_field_type_1_is_repeated : _GEN_5825; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5827 = _GEN_11169 & _GEN_10646 ? field_stack_8_field_type_2_is_repeated : _GEN_5826; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5828 = _GEN_11169 & _GEN_10648 ? field_stack_8_field_type_3_is_repeated : _GEN_5827; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5829 = _GEN_11169 & _GEN_10650 ? field_stack_8_field_type_4_is_repeated : _GEN_5828; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5830 = _GEN_11169 & _GEN_10652 ? field_stack_8_field_type_5_is_repeated : _GEN_5829; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5831 = _GEN_11169 & _GEN_10654 ? field_stack_8_field_type_6_is_repeated : _GEN_5830; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5832 = _GEN_11169 & _GEN_10656 ? field_stack_8_field_type_7_is_repeated : _GEN_5831; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5833 = _GEN_11169 & _GEN_10658 ? field_stack_8_field_type_8_is_repeated : _GEN_5832; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5834 = _GEN_11169 & _GEN_10660 ? field_stack_8_field_type_9_is_repeated : _GEN_5833; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5835 = _GEN_11169 & _GEN_10662 ? field_stack_8_field_type_10_is_repeated : _GEN_5834; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5836 = _GEN_11169 & _GEN_10664 ? field_stack_8_field_type_11_is_repeated : _GEN_5835; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5837 = _GEN_11169 & _GEN_10666 ? field_stack_8_field_type_12_is_repeated : _GEN_5836; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5838 = _GEN_11169 & _GEN_10668 ? field_stack_8_field_type_13_is_repeated : _GEN_5837; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5839 = _GEN_11169 & _GEN_10670 ? field_stack_8_field_type_14_is_repeated : _GEN_5838; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5840 = _GEN_11169 & _GEN_10672 ? field_stack_8_field_type_15_is_repeated : _GEN_5839; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5841 = _GEN_11169 & _GEN_10674 ? field_stack_8_field_type_16_is_repeated : _GEN_5840; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5842 = _GEN_11169 & _GEN_10676 ? field_stack_8_field_type_17_is_repeated : _GEN_5841; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5843 = _GEN_11169 & _GEN_10678 ? field_stack_8_field_type_18_is_repeated : _GEN_5842; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5844 = _GEN_11169 & _GEN_10680 ? field_stack_8_field_type_19_is_repeated : _GEN_5843; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5845 = _GEN_11169 & _GEN_10682 ? field_stack_8_field_type_20_is_repeated : _GEN_5844; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5846 = _GEN_11169 & _GEN_10684 ? field_stack_8_field_type_21_is_repeated : _GEN_5845; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5847 = _GEN_11169 & _GEN_10686 ? field_stack_8_field_type_22_is_repeated : _GEN_5846; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5848 = _GEN_11169 & _GEN_10688 ? field_stack_8_field_type_23_is_repeated : _GEN_5847; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5849 = _GEN_11169 & _GEN_10690 ? field_stack_8_field_type_24_is_repeated : _GEN_5848; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5850 = _GEN_11169 & _GEN_10692 ? field_stack_8_field_type_25_is_repeated : _GEN_5849; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5851 = _GEN_11169 & _GEN_10694 ? field_stack_8_field_type_26_is_repeated : _GEN_5850; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5852 = _GEN_11169 & _GEN_10696 ? field_stack_8_field_type_27_is_repeated : _GEN_5851; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5853 = _GEN_11169 & _GEN_10698 ? field_stack_8_field_type_28_is_repeated : _GEN_5852; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5854 = _GEN_11169 & _GEN_10700 ? field_stack_8_field_type_29_is_repeated : _GEN_5853; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5855 = _GEN_11169 & _GEN_10702 ? field_stack_8_field_type_30_is_repeated : _GEN_5854; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5856 = _GEN_11169 & _GEN_10704 ? field_stack_8_field_type_31_is_repeated : _GEN_5855; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5857 = _GEN_11169 & _GEN_10706 ? field_stack_8_field_type_32_is_repeated : _GEN_5856; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5858 = _GEN_11235 & _GEN_10708 ? field_stack_9_field_type_0_is_repeated : _GEN_5857; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5859 = _GEN_11235 & _GEN_10644 ? field_stack_9_field_type_1_is_repeated : _GEN_5858; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5860 = _GEN_11235 & _GEN_10646 ? field_stack_9_field_type_2_is_repeated : _GEN_5859; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5861 = _GEN_11235 & _GEN_10648 ? field_stack_9_field_type_3_is_repeated : _GEN_5860; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5862 = _GEN_11235 & _GEN_10650 ? field_stack_9_field_type_4_is_repeated : _GEN_5861; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5863 = _GEN_11235 & _GEN_10652 ? field_stack_9_field_type_5_is_repeated : _GEN_5862; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5864 = _GEN_11235 & _GEN_10654 ? field_stack_9_field_type_6_is_repeated : _GEN_5863; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5865 = _GEN_11235 & _GEN_10656 ? field_stack_9_field_type_7_is_repeated : _GEN_5864; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5866 = _GEN_11235 & _GEN_10658 ? field_stack_9_field_type_8_is_repeated : _GEN_5865; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5867 = _GEN_11235 & _GEN_10660 ? field_stack_9_field_type_9_is_repeated : _GEN_5866; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5868 = _GEN_11235 & _GEN_10662 ? field_stack_9_field_type_10_is_repeated : _GEN_5867; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5869 = _GEN_11235 & _GEN_10664 ? field_stack_9_field_type_11_is_repeated : _GEN_5868; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5870 = _GEN_11235 & _GEN_10666 ? field_stack_9_field_type_12_is_repeated : _GEN_5869; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5871 = _GEN_11235 & _GEN_10668 ? field_stack_9_field_type_13_is_repeated : _GEN_5870; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5872 = _GEN_11235 & _GEN_10670 ? field_stack_9_field_type_14_is_repeated : _GEN_5871; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5873 = _GEN_11235 & _GEN_10672 ? field_stack_9_field_type_15_is_repeated : _GEN_5872; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5874 = _GEN_11235 & _GEN_10674 ? field_stack_9_field_type_16_is_repeated : _GEN_5873; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5875 = _GEN_11235 & _GEN_10676 ? field_stack_9_field_type_17_is_repeated : _GEN_5874; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5876 = _GEN_11235 & _GEN_10678 ? field_stack_9_field_type_18_is_repeated : _GEN_5875; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5877 = _GEN_11235 & _GEN_10680 ? field_stack_9_field_type_19_is_repeated : _GEN_5876; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5878 = _GEN_11235 & _GEN_10682 ? field_stack_9_field_type_20_is_repeated : _GEN_5877; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5879 = _GEN_11235 & _GEN_10684 ? field_stack_9_field_type_21_is_repeated : _GEN_5878; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5880 = _GEN_11235 & _GEN_10686 ? field_stack_9_field_type_22_is_repeated : _GEN_5879; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5881 = _GEN_11235 & _GEN_10688 ? field_stack_9_field_type_23_is_repeated : _GEN_5880; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5882 = _GEN_11235 & _GEN_10690 ? field_stack_9_field_type_24_is_repeated : _GEN_5881; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5883 = _GEN_11235 & _GEN_10692 ? field_stack_9_field_type_25_is_repeated : _GEN_5882; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5884 = _GEN_11235 & _GEN_10694 ? field_stack_9_field_type_26_is_repeated : _GEN_5883; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5885 = _GEN_11235 & _GEN_10696 ? field_stack_9_field_type_27_is_repeated : _GEN_5884; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5886 = _GEN_11235 & _GEN_10698 ? field_stack_9_field_type_28_is_repeated : _GEN_5885; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5887 = _GEN_11235 & _GEN_10700 ? field_stack_9_field_type_29_is_repeated : _GEN_5886; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5888 = _GEN_11235 & _GEN_10702 ? field_stack_9_field_type_30_is_repeated : _GEN_5887; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5889 = _GEN_11235 & _GEN_10704 ? field_stack_9_field_type_31_is_repeated : _GEN_5888; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5890 = _GEN_11235 & _GEN_10706 ? field_stack_9_field_type_32_is_repeated : _GEN_5889; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5891 = _GEN_11301 & _GEN_10708 ? field_stack_10_field_type_0_is_repeated : _GEN_5890; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5892 = _GEN_11301 & _GEN_10644 ? field_stack_10_field_type_1_is_repeated : _GEN_5891; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5893 = _GEN_11301 & _GEN_10646 ? field_stack_10_field_type_2_is_repeated : _GEN_5892; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5894 = _GEN_11301 & _GEN_10648 ? field_stack_10_field_type_3_is_repeated : _GEN_5893; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5895 = _GEN_11301 & _GEN_10650 ? field_stack_10_field_type_4_is_repeated : _GEN_5894; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5896 = _GEN_11301 & _GEN_10652 ? field_stack_10_field_type_5_is_repeated : _GEN_5895; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5897 = _GEN_11301 & _GEN_10654 ? field_stack_10_field_type_6_is_repeated : _GEN_5896; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5898 = _GEN_11301 & _GEN_10656 ? field_stack_10_field_type_7_is_repeated : _GEN_5897; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5899 = _GEN_11301 & _GEN_10658 ? field_stack_10_field_type_8_is_repeated : _GEN_5898; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5900 = _GEN_11301 & _GEN_10660 ? field_stack_10_field_type_9_is_repeated : _GEN_5899; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5901 = _GEN_11301 & _GEN_10662 ? field_stack_10_field_type_10_is_repeated : _GEN_5900; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5902 = _GEN_11301 & _GEN_10664 ? field_stack_10_field_type_11_is_repeated : _GEN_5901; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5903 = _GEN_11301 & _GEN_10666 ? field_stack_10_field_type_12_is_repeated : _GEN_5902; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5904 = _GEN_11301 & _GEN_10668 ? field_stack_10_field_type_13_is_repeated : _GEN_5903; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5905 = _GEN_11301 & _GEN_10670 ? field_stack_10_field_type_14_is_repeated : _GEN_5904; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5906 = _GEN_11301 & _GEN_10672 ? field_stack_10_field_type_15_is_repeated : _GEN_5905; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5907 = _GEN_11301 & _GEN_10674 ? field_stack_10_field_type_16_is_repeated : _GEN_5906; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5908 = _GEN_11301 & _GEN_10676 ? field_stack_10_field_type_17_is_repeated : _GEN_5907; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5909 = _GEN_11301 & _GEN_10678 ? field_stack_10_field_type_18_is_repeated : _GEN_5908; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5910 = _GEN_11301 & _GEN_10680 ? field_stack_10_field_type_19_is_repeated : _GEN_5909; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5911 = _GEN_11301 & _GEN_10682 ? field_stack_10_field_type_20_is_repeated : _GEN_5910; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5912 = _GEN_11301 & _GEN_10684 ? field_stack_10_field_type_21_is_repeated : _GEN_5911; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5913 = _GEN_11301 & _GEN_10686 ? field_stack_10_field_type_22_is_repeated : _GEN_5912; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5914 = _GEN_11301 & _GEN_10688 ? field_stack_10_field_type_23_is_repeated : _GEN_5913; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5915 = _GEN_11301 & _GEN_10690 ? field_stack_10_field_type_24_is_repeated : _GEN_5914; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5916 = _GEN_11301 & _GEN_10692 ? field_stack_10_field_type_25_is_repeated : _GEN_5915; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5917 = _GEN_11301 & _GEN_10694 ? field_stack_10_field_type_26_is_repeated : _GEN_5916; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5918 = _GEN_11301 & _GEN_10696 ? field_stack_10_field_type_27_is_repeated : _GEN_5917; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5919 = _GEN_11301 & _GEN_10698 ? field_stack_10_field_type_28_is_repeated : _GEN_5918; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5920 = _GEN_11301 & _GEN_10700 ? field_stack_10_field_type_29_is_repeated : _GEN_5919; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5921 = _GEN_11301 & _GEN_10702 ? field_stack_10_field_type_30_is_repeated : _GEN_5920; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5922 = _GEN_11301 & _GEN_10704 ? field_stack_10_field_type_31_is_repeated : _GEN_5921; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5923 = _GEN_11301 & _GEN_10706 ? field_stack_10_field_type_32_is_repeated : _GEN_5922; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5924 = _GEN_11367 & _GEN_10708 ? field_stack_11_field_type_0_is_repeated : _GEN_5923; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5925 = _GEN_11367 & _GEN_10644 ? field_stack_11_field_type_1_is_repeated : _GEN_5924; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5926 = _GEN_11367 & _GEN_10646 ? field_stack_11_field_type_2_is_repeated : _GEN_5925; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5927 = _GEN_11367 & _GEN_10648 ? field_stack_11_field_type_3_is_repeated : _GEN_5926; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5928 = _GEN_11367 & _GEN_10650 ? field_stack_11_field_type_4_is_repeated : _GEN_5927; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5929 = _GEN_11367 & _GEN_10652 ? field_stack_11_field_type_5_is_repeated : _GEN_5928; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5930 = _GEN_11367 & _GEN_10654 ? field_stack_11_field_type_6_is_repeated : _GEN_5929; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5931 = _GEN_11367 & _GEN_10656 ? field_stack_11_field_type_7_is_repeated : _GEN_5930; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5932 = _GEN_11367 & _GEN_10658 ? field_stack_11_field_type_8_is_repeated : _GEN_5931; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5933 = _GEN_11367 & _GEN_10660 ? field_stack_11_field_type_9_is_repeated : _GEN_5932; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5934 = _GEN_11367 & _GEN_10662 ? field_stack_11_field_type_10_is_repeated : _GEN_5933; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5935 = _GEN_11367 & _GEN_10664 ? field_stack_11_field_type_11_is_repeated : _GEN_5934; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5936 = _GEN_11367 & _GEN_10666 ? field_stack_11_field_type_12_is_repeated : _GEN_5935; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5937 = _GEN_11367 & _GEN_10668 ? field_stack_11_field_type_13_is_repeated : _GEN_5936; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5938 = _GEN_11367 & _GEN_10670 ? field_stack_11_field_type_14_is_repeated : _GEN_5937; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5939 = _GEN_11367 & _GEN_10672 ? field_stack_11_field_type_15_is_repeated : _GEN_5938; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5940 = _GEN_11367 & _GEN_10674 ? field_stack_11_field_type_16_is_repeated : _GEN_5939; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5941 = _GEN_11367 & _GEN_10676 ? field_stack_11_field_type_17_is_repeated : _GEN_5940; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5942 = _GEN_11367 & _GEN_10678 ? field_stack_11_field_type_18_is_repeated : _GEN_5941; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5943 = _GEN_11367 & _GEN_10680 ? field_stack_11_field_type_19_is_repeated : _GEN_5942; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5944 = _GEN_11367 & _GEN_10682 ? field_stack_11_field_type_20_is_repeated : _GEN_5943; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5945 = _GEN_11367 & _GEN_10684 ? field_stack_11_field_type_21_is_repeated : _GEN_5944; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5946 = _GEN_11367 & _GEN_10686 ? field_stack_11_field_type_22_is_repeated : _GEN_5945; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5947 = _GEN_11367 & _GEN_10688 ? field_stack_11_field_type_23_is_repeated : _GEN_5946; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5948 = _GEN_11367 & _GEN_10690 ? field_stack_11_field_type_24_is_repeated : _GEN_5947; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5949 = _GEN_11367 & _GEN_10692 ? field_stack_11_field_type_25_is_repeated : _GEN_5948; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5950 = _GEN_11367 & _GEN_10694 ? field_stack_11_field_type_26_is_repeated : _GEN_5949; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5951 = _GEN_11367 & _GEN_10696 ? field_stack_11_field_type_27_is_repeated : _GEN_5950; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5952 = _GEN_11367 & _GEN_10698 ? field_stack_11_field_type_28_is_repeated : _GEN_5951; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5953 = _GEN_11367 & _GEN_10700 ? field_stack_11_field_type_29_is_repeated : _GEN_5952; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5954 = _GEN_11367 & _GEN_10702 ? field_stack_11_field_type_30_is_repeated : _GEN_5953; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5955 = _GEN_11367 & _GEN_10704 ? field_stack_11_field_type_31_is_repeated : _GEN_5954; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5956 = _GEN_11367 & _GEN_10706 ? field_stack_11_field_type_32_is_repeated : _GEN_5955; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5957 = _GEN_11433 & _GEN_10708 ? field_stack_12_field_type_0_is_repeated : _GEN_5956; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5958 = _GEN_11433 & _GEN_10644 ? field_stack_12_field_type_1_is_repeated : _GEN_5957; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5959 = _GEN_11433 & _GEN_10646 ? field_stack_12_field_type_2_is_repeated : _GEN_5958; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5960 = _GEN_11433 & _GEN_10648 ? field_stack_12_field_type_3_is_repeated : _GEN_5959; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5961 = _GEN_11433 & _GEN_10650 ? field_stack_12_field_type_4_is_repeated : _GEN_5960; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5962 = _GEN_11433 & _GEN_10652 ? field_stack_12_field_type_5_is_repeated : _GEN_5961; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5963 = _GEN_11433 & _GEN_10654 ? field_stack_12_field_type_6_is_repeated : _GEN_5962; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5964 = _GEN_11433 & _GEN_10656 ? field_stack_12_field_type_7_is_repeated : _GEN_5963; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5965 = _GEN_11433 & _GEN_10658 ? field_stack_12_field_type_8_is_repeated : _GEN_5964; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5966 = _GEN_11433 & _GEN_10660 ? field_stack_12_field_type_9_is_repeated : _GEN_5965; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5967 = _GEN_11433 & _GEN_10662 ? field_stack_12_field_type_10_is_repeated : _GEN_5966; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5968 = _GEN_11433 & _GEN_10664 ? field_stack_12_field_type_11_is_repeated : _GEN_5967; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5969 = _GEN_11433 & _GEN_10666 ? field_stack_12_field_type_12_is_repeated : _GEN_5968; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5970 = _GEN_11433 & _GEN_10668 ? field_stack_12_field_type_13_is_repeated : _GEN_5969; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5971 = _GEN_11433 & _GEN_10670 ? field_stack_12_field_type_14_is_repeated : _GEN_5970; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5972 = _GEN_11433 & _GEN_10672 ? field_stack_12_field_type_15_is_repeated : _GEN_5971; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5973 = _GEN_11433 & _GEN_10674 ? field_stack_12_field_type_16_is_repeated : _GEN_5972; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5974 = _GEN_11433 & _GEN_10676 ? field_stack_12_field_type_17_is_repeated : _GEN_5973; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5975 = _GEN_11433 & _GEN_10678 ? field_stack_12_field_type_18_is_repeated : _GEN_5974; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5976 = _GEN_11433 & _GEN_10680 ? field_stack_12_field_type_19_is_repeated : _GEN_5975; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5977 = _GEN_11433 & _GEN_10682 ? field_stack_12_field_type_20_is_repeated : _GEN_5976; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5978 = _GEN_11433 & _GEN_10684 ? field_stack_12_field_type_21_is_repeated : _GEN_5977; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5979 = _GEN_11433 & _GEN_10686 ? field_stack_12_field_type_22_is_repeated : _GEN_5978; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5980 = _GEN_11433 & _GEN_10688 ? field_stack_12_field_type_23_is_repeated : _GEN_5979; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5981 = _GEN_11433 & _GEN_10690 ? field_stack_12_field_type_24_is_repeated : _GEN_5980; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5982 = _GEN_11433 & _GEN_10692 ? field_stack_12_field_type_25_is_repeated : _GEN_5981; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5983 = _GEN_11433 & _GEN_10694 ? field_stack_12_field_type_26_is_repeated : _GEN_5982; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5984 = _GEN_11433 & _GEN_10696 ? field_stack_12_field_type_27_is_repeated : _GEN_5983; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5985 = _GEN_11433 & _GEN_10698 ? field_stack_12_field_type_28_is_repeated : _GEN_5984; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5986 = _GEN_11433 & _GEN_10700 ? field_stack_12_field_type_29_is_repeated : _GEN_5985; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5987 = _GEN_11433 & _GEN_10702 ? field_stack_12_field_type_30_is_repeated : _GEN_5986; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5988 = _GEN_11433 & _GEN_10704 ? field_stack_12_field_type_31_is_repeated : _GEN_5987; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5989 = _GEN_11433 & _GEN_10706 ? field_stack_12_field_type_32_is_repeated : _GEN_5988; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5990 = _GEN_11499 & _GEN_10708 ? field_stack_13_field_type_0_is_repeated : _GEN_5989; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5991 = _GEN_11499 & _GEN_10644 ? field_stack_13_field_type_1_is_repeated : _GEN_5990; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5992 = _GEN_11499 & _GEN_10646 ? field_stack_13_field_type_2_is_repeated : _GEN_5991; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5993 = _GEN_11499 & _GEN_10648 ? field_stack_13_field_type_3_is_repeated : _GEN_5992; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5994 = _GEN_11499 & _GEN_10650 ? field_stack_13_field_type_4_is_repeated : _GEN_5993; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5995 = _GEN_11499 & _GEN_10652 ? field_stack_13_field_type_5_is_repeated : _GEN_5994; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5996 = _GEN_11499 & _GEN_10654 ? field_stack_13_field_type_6_is_repeated : _GEN_5995; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5997 = _GEN_11499 & _GEN_10656 ? field_stack_13_field_type_7_is_repeated : _GEN_5996; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5998 = _GEN_11499 & _GEN_10658 ? field_stack_13_field_type_8_is_repeated : _GEN_5997; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_5999 = _GEN_11499 & _GEN_10660 ? field_stack_13_field_type_9_is_repeated : _GEN_5998; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_6000 = _GEN_11499 & _GEN_10662 ? field_stack_13_field_type_10_is_repeated : _GEN_5999; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_6001 = _GEN_11499 & _GEN_10664 ? field_stack_13_field_type_11_is_repeated : _GEN_6000; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_6002 = _GEN_11499 & _GEN_10666 ? field_stack_13_field_type_12_is_repeated : _GEN_6001; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_6003 = _GEN_11499 & _GEN_10668 ? field_stack_13_field_type_13_is_repeated : _GEN_6002; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_6004 = _GEN_11499 & _GEN_10670 ? field_stack_13_field_type_14_is_repeated : _GEN_6003; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_6005 = _GEN_11499 & _GEN_10672 ? field_stack_13_field_type_15_is_repeated : _GEN_6004; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_6006 = _GEN_11499 & _GEN_10674 ? field_stack_13_field_type_16_is_repeated : _GEN_6005; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_6007 = _GEN_11499 & _GEN_10676 ? field_stack_13_field_type_17_is_repeated : _GEN_6006; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_6008 = _GEN_11499 & _GEN_10678 ? field_stack_13_field_type_18_is_repeated : _GEN_6007; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_6009 = _GEN_11499 & _GEN_10680 ? field_stack_13_field_type_19_is_repeated : _GEN_6008; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_6010 = _GEN_11499 & _GEN_10682 ? field_stack_13_field_type_20_is_repeated : _GEN_6009; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_6011 = _GEN_11499 & _GEN_10684 ? field_stack_13_field_type_21_is_repeated : _GEN_6010; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_6012 = _GEN_11499 & _GEN_10686 ? field_stack_13_field_type_22_is_repeated : _GEN_6011; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_6013 = _GEN_11499 & _GEN_10688 ? field_stack_13_field_type_23_is_repeated : _GEN_6012; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_6014 = _GEN_11499 & _GEN_10690 ? field_stack_13_field_type_24_is_repeated : _GEN_6013; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_6015 = _GEN_11499 & _GEN_10692 ? field_stack_13_field_type_25_is_repeated : _GEN_6014; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_6016 = _GEN_11499 & _GEN_10694 ? field_stack_13_field_type_26_is_repeated : _GEN_6015; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_6017 = _GEN_11499 & _GEN_10696 ? field_stack_13_field_type_27_is_repeated : _GEN_6016; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_6018 = _GEN_11499 & _GEN_10698 ? field_stack_13_field_type_28_is_repeated : _GEN_6017; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_6019 = _GEN_11499 & _GEN_10700 ? field_stack_13_field_type_29_is_repeated : _GEN_6018; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_6020 = _GEN_11499 & _GEN_10702 ? field_stack_13_field_type_30_is_repeated : _GEN_6019; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_6021 = _GEN_11499 & _GEN_10704 ? field_stack_13_field_type_31_is_repeated : _GEN_6020; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_6022 = _GEN_11499 & _GEN_10706 ? field_stack_13_field_type_32_is_repeated : _GEN_6021; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_6023 = _GEN_11565 & _GEN_10708 ? field_stack_14_field_type_0_is_repeated : _GEN_6022; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_6024 = _GEN_11565 & _GEN_10644 ? field_stack_14_field_type_1_is_repeated : _GEN_6023; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_6025 = _GEN_11565 & _GEN_10646 ? field_stack_14_field_type_2_is_repeated : _GEN_6024; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_6026 = _GEN_11565 & _GEN_10648 ? field_stack_14_field_type_3_is_repeated : _GEN_6025; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_6027 = _GEN_11565 & _GEN_10650 ? field_stack_14_field_type_4_is_repeated : _GEN_6026; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_6028 = _GEN_11565 & _GEN_10652 ? field_stack_14_field_type_5_is_repeated : _GEN_6027; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_6029 = _GEN_11565 & _GEN_10654 ? field_stack_14_field_type_6_is_repeated : _GEN_6028; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_6030 = _GEN_11565 & _GEN_10656 ? field_stack_14_field_type_7_is_repeated : _GEN_6029; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_6031 = _GEN_11565 & _GEN_10658 ? field_stack_14_field_type_8_is_repeated : _GEN_6030; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_6032 = _GEN_11565 & _GEN_10660 ? field_stack_14_field_type_9_is_repeated : _GEN_6031; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_6033 = _GEN_11565 & _GEN_10662 ? field_stack_14_field_type_10_is_repeated : _GEN_6032; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_6034 = _GEN_11565 & _GEN_10664 ? field_stack_14_field_type_11_is_repeated : _GEN_6033; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_6035 = _GEN_11565 & _GEN_10666 ? field_stack_14_field_type_12_is_repeated : _GEN_6034; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_6036 = _GEN_11565 & _GEN_10668 ? field_stack_14_field_type_13_is_repeated : _GEN_6035; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_6037 = _GEN_11565 & _GEN_10670 ? field_stack_14_field_type_14_is_repeated : _GEN_6036; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_6038 = _GEN_11565 & _GEN_10672 ? field_stack_14_field_type_15_is_repeated : _GEN_6037; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_6039 = _GEN_11565 & _GEN_10674 ? field_stack_14_field_type_16_is_repeated : _GEN_6038; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_6040 = _GEN_11565 & _GEN_10676 ? field_stack_14_field_type_17_is_repeated : _GEN_6039; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_6041 = _GEN_11565 & _GEN_10678 ? field_stack_14_field_type_18_is_repeated : _GEN_6040; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_6042 = _GEN_11565 & _GEN_10680 ? field_stack_14_field_type_19_is_repeated : _GEN_6041; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_6043 = _GEN_11565 & _GEN_10682 ? field_stack_14_field_type_20_is_repeated : _GEN_6042; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_6044 = _GEN_11565 & _GEN_10684 ? field_stack_14_field_type_21_is_repeated : _GEN_6043; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_6045 = _GEN_11565 & _GEN_10686 ? field_stack_14_field_type_22_is_repeated : _GEN_6044; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_6046 = _GEN_11565 & _GEN_10688 ? field_stack_14_field_type_23_is_repeated : _GEN_6045; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_6047 = _GEN_11565 & _GEN_10690 ? field_stack_14_field_type_24_is_repeated : _GEN_6046; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_6048 = _GEN_11565 & _GEN_10692 ? field_stack_14_field_type_25_is_repeated : _GEN_6047; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_6049 = _GEN_11565 & _GEN_10694 ? field_stack_14_field_type_26_is_repeated : _GEN_6048; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_6050 = _GEN_11565 & _GEN_10696 ? field_stack_14_field_type_27_is_repeated : _GEN_6049; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_6051 = _GEN_11565 & _GEN_10698 ? field_stack_14_field_type_28_is_repeated : _GEN_6050; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_6052 = _GEN_11565 & _GEN_10700 ? field_stack_14_field_type_29_is_repeated : _GEN_6051; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_6053 = _GEN_11565 & _GEN_10702 ? field_stack_14_field_type_30_is_repeated : _GEN_6052; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_6054 = _GEN_11565 & _GEN_10704 ? field_stack_14_field_type_31_is_repeated : _GEN_6053; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire  _GEN_6055 = _GEN_11565 & _GEN_10706 ? field_stack_14_field_type_32_is_repeated : _GEN_6054; // @[Serializerhw.scala 140:45 Serializerhw.scala 140:45]
  wire [4:0] _GEN_6056 = _GEN_4570 == 5'h0 ? 5'h13 : 5'h12; // @[Serializerhw.scala 136:98 Serializerhw.scala 137:45 Serializerhw.scala 141:45]
  wire [5:0] _GEN_6057 = _GEN_4570 == 5'h0 ? _current_field_num_T_1 : current_field_num; // @[Serializerhw.scala 136:98 Serializerhw.scala 138:45 Serializerhw.scala 73:36]
  wire [15:0] _GEN_6059 = _GEN_4570 == 5'h0 ? c_sub_metadata_sub_class_id : _GEN_5560; // @[Serializerhw.scala 136:98 Serializerhw.scala 74:33 Serializerhw.scala 140:45]
  wire [4:0] _GEN_6060 = _GEN_4570 == 5'h0 ? c_sub_metadata_field_type : _GEN_4570; // @[Serializerhw.scala 136:98 Serializerhw.scala 74:33 Serializerhw.scala 140:45]
  wire  _GEN_6061 = _GEN_4570 == 5'h0 ? c_sub_metadata_is_repeated : _GEN_6055; // @[Serializerhw.scala 136:98 Serializerhw.scala 74:33 Serializerhw.scala 140:45]
  wire [4:0] _GEN_6062 = current_field_num == 6'h0 ? _GEN_4075 : _GEN_6056; // @[Serializerhw.scala 130:44]
  wire [5:0] _GEN_6063 = current_field_num == 6'h0 ? current_field_num : _GEN_6057; // @[Serializerhw.scala 130:44 Serializerhw.scala 73:36]
  wire [15:0] _GEN_6065 = current_field_num == 6'h0 ? c_sub_metadata_sub_class_id : _GEN_6059; // @[Serializerhw.scala 130:44 Serializerhw.scala 74:33]
  wire [4:0] _GEN_6066 = current_field_num == 6'h0 ? c_sub_metadata_field_type : _GEN_6060; // @[Serializerhw.scala 130:44 Serializerhw.scala 74:33]
  wire  _GEN_6067 = current_field_num == 6'h0 ? c_sub_metadata_is_repeated : _GEN_6061; // @[Serializerhw.scala 130:44 Serializerhw.scala 74:33]
  wire  _T_14 = 5'h12 == state; // @[Conditional.scala 37:30]
  wire [2:0] _GEN_6069 = 5'h1 == c_sub_metadata_field_type ? 3'h1 : 3'h0; // @[Serializerhw.scala 147:84 Serializerhw.scala 147:84]
  wire [2:0] _GEN_6070 = 5'h2 == c_sub_metadata_field_type ? 3'h5 : _GEN_6069; // @[Serializerhw.scala 147:84 Serializerhw.scala 147:84]
  wire [2:0] _GEN_6071 = 5'h3 == c_sub_metadata_field_type ? 3'h0 : _GEN_6070; // @[Serializerhw.scala 147:84 Serializerhw.scala 147:84]
  wire [2:0] _GEN_6072 = 5'h4 == c_sub_metadata_field_type ? 3'h0 : _GEN_6071; // @[Serializerhw.scala 147:84 Serializerhw.scala 147:84]
  wire [2:0] _GEN_6073 = 5'h5 == c_sub_metadata_field_type ? 3'h0 : _GEN_6072; // @[Serializerhw.scala 147:84 Serializerhw.scala 147:84]
  wire [2:0] _GEN_6074 = 5'h6 == c_sub_metadata_field_type ? 3'h1 : _GEN_6073; // @[Serializerhw.scala 147:84 Serializerhw.scala 147:84]
  wire [2:0] _GEN_6075 = 5'h7 == c_sub_metadata_field_type ? 3'h5 : _GEN_6074; // @[Serializerhw.scala 147:84 Serializerhw.scala 147:84]
  wire [2:0] _GEN_6076 = 5'h8 == c_sub_metadata_field_type ? 3'h0 : _GEN_6075; // @[Serializerhw.scala 147:84 Serializerhw.scala 147:84]
  wire [2:0] _GEN_6077 = 5'h9 == c_sub_metadata_field_type ? 3'h2 : _GEN_6076; // @[Serializerhw.scala 147:84 Serializerhw.scala 147:84]
  wire [2:0] _GEN_6078 = 5'ha == c_sub_metadata_field_type ? 3'h3 : _GEN_6077; // @[Serializerhw.scala 147:84 Serializerhw.scala 147:84]
  wire [2:0] _GEN_6079 = 5'hb == c_sub_metadata_field_type ? 3'h2 : _GEN_6078; // @[Serializerhw.scala 147:84 Serializerhw.scala 147:84]
  wire [2:0] _GEN_6080 = 5'hc == c_sub_metadata_field_type ? 3'h2 : _GEN_6079; // @[Serializerhw.scala 147:84 Serializerhw.scala 147:84]
  wire [2:0] _GEN_6081 = 5'hd == c_sub_metadata_field_type ? 3'h0 : _GEN_6080; // @[Serializerhw.scala 147:84 Serializerhw.scala 147:84]
  wire [2:0] _GEN_6082 = 5'he == c_sub_metadata_field_type ? 3'h0 : _GEN_6081; // @[Serializerhw.scala 147:84 Serializerhw.scala 147:84]
  wire [2:0] _GEN_6083 = 5'hf == c_sub_metadata_field_type ? 3'h5 : _GEN_6082; // @[Serializerhw.scala 147:84 Serializerhw.scala 147:84]
  wire [2:0] _GEN_6084 = 5'h10 == c_sub_metadata_field_type ? 3'h1 : _GEN_6083; // @[Serializerhw.scala 147:84 Serializerhw.scala 147:84]
  wire [2:0] _GEN_6085 = 5'h11 == c_sub_metadata_field_type ? 3'h0 : _GEN_6084; // @[Serializerhw.scala 147:84 Serializerhw.scala 147:84]
  wire [2:0] _GEN_6086 = 5'h12 == c_sub_metadata_field_type ? 3'h0 : _GEN_6085; // @[Serializerhw.scala 147:84 Serializerhw.scala 147:84]
  wire [4:0] _GEN_6125 = _GEN_6086 == 3'h5 ? 5'h5 : 5'h2; // @[Serializerhw.scala 151:121 Serializerhw.scala 152:41 Serializerhw.scala 154:41]
  wire [4:0] _GEN_6126 = _GEN_6086 == 3'h1 ? 5'h1 : _GEN_6125; // @[Serializerhw.scala 149:121 Serializerhw.scala 150:41]
  wire [4:0] _GEN_6127 = _GEN_6086 == 3'h0 ? 5'h0 : _GEN_6126; // @[Serializerhw.scala 147:116 Serializerhw.scala 148:41]
  wire [15:0] _GEN_6188 = c_sub_metadata_is_repeated ? c_sub_metadata_sub_class_id : 16'h0; // @[Serializerhw.scala 145:45 Serializerhw.scala 146:41 Serializerhw.scala 158:41]
  wire [4:0] _GEN_6189 = c_sub_metadata_is_repeated ? _GEN_6127 : _GEN_6127; // @[Serializerhw.scala 145:45]
  wire  _T_21 = 5'h0 == state; // @[Conditional.scala 37:30]
  wire  _T_22 = repeat_num == 8'h0; // @[Serializerhw.scala 171:29]
  wire  _T_23 = repeat_num == 8'h1; // @[Serializerhw.scala 174:35]
  wire [7:0] _repeat_num_T_1 = repeat_num - 8'h1; // @[Serializerhw.scala 178:67]
  wire [4:0] _GEN_6190 = repeat_num == 8'h1 ? 5'hc : 5'h0; // @[Serializerhw.scala 174:43 Serializerhw.scala 175:45 Serializerhw.scala 177:53]
  wire [7:0] _GEN_6191 = repeat_num == 8'h1 ? repeat_num : _repeat_num_T_1; // @[Serializerhw.scala 174:43 Serializerhw.scala 75:29 Serializerhw.scala 178:53]
  wire [4:0] _GEN_6192 = repeat_num == 8'h0 ? 5'h13 : _GEN_6190; // @[Serializerhw.scala 171:37 Serializerhw.scala 172:45]
  wire [5:0] _GEN_6193 = repeat_num == 8'h0 ? _current_field_num_T_1 : current_field_num; // @[Serializerhw.scala 171:37 Serializerhw.scala 173:45 Serializerhw.scala 73:36]
  wire [7:0] _GEN_6194 = repeat_num == 8'h0 ? repeat_num : _GEN_6191; // @[Serializerhw.scala 171:37 Serializerhw.scala 75:29]
  wire  _T_24 = 5'h5 == state; // @[Conditional.scala 37:30]
  wire [4:0] _GEN_6195 = _T_23 ? 5'hc : 5'h5; // @[Serializerhw.scala 185:43 Serializerhw.scala 186:45 Serializerhw.scala 188:53]
  wire [4:0] _GEN_6197 = _T_22 ? 5'h13 : _GEN_6195; // @[Serializerhw.scala 182:37 Serializerhw.scala 183:45]
  wire  _T_27 = 5'h1 == state; // @[Conditional.scala 37:30]
  wire [4:0] _GEN_6200 = _T_23 ? 5'hc : state; // @[Serializerhw.scala 196:43 Serializerhw.scala 197:45 Serializerhw.scala 86:46]
  wire [4:0] _GEN_6202 = _T_22 ? 5'h13 : _GEN_6200; // @[Serializerhw.scala 193:37 Serializerhw.scala 194:45]
  wire  _T_30 = 5'h2 == state; // @[Conditional.scala 37:30]
  wire  _T_31 = c_sub_metadata_field_type == 5'hb; // @[Serializerhw.scala 203:46]
  wire [3:0] _stack_num_T_1 = stack_num + 4'h1; // @[Serializerhw.scala 206:70]
  wire [5:0] _GEN_6205 = 4'h0 == stack_num ? current_field_num : field_num_0; // @[Serializerhw.scala 207:57 Serializerhw.scala 207:57 Serializerhw.scala 70:28]
  wire [5:0] _GEN_6206 = 4'h1 == stack_num ? current_field_num : field_num_1; // @[Serializerhw.scala 207:57 Serializerhw.scala 207:57 Serializerhw.scala 70:28]
  wire [5:0] _GEN_6207 = 4'h2 == stack_num ? current_field_num : field_num_2; // @[Serializerhw.scala 207:57 Serializerhw.scala 207:57 Serializerhw.scala 70:28]
  wire [5:0] _GEN_6208 = 4'h3 == stack_num ? current_field_num : field_num_3; // @[Serializerhw.scala 207:57 Serializerhw.scala 207:57 Serializerhw.scala 70:28]
  wire [5:0] _GEN_6209 = 4'h4 == stack_num ? current_field_num : field_num_4; // @[Serializerhw.scala 207:57 Serializerhw.scala 207:57 Serializerhw.scala 70:28]
  wire [5:0] _GEN_6210 = 4'h5 == stack_num ? current_field_num : field_num_5; // @[Serializerhw.scala 207:57 Serializerhw.scala 207:57 Serializerhw.scala 70:28]
  wire [5:0] _GEN_6211 = 4'h6 == stack_num ? current_field_num : field_num_6; // @[Serializerhw.scala 207:57 Serializerhw.scala 207:57 Serializerhw.scala 70:28]
  wire [5:0] _GEN_6212 = 4'h7 == stack_num ? current_field_num : field_num_7; // @[Serializerhw.scala 207:57 Serializerhw.scala 207:57 Serializerhw.scala 70:28]
  wire [5:0] _GEN_6213 = 4'h8 == stack_num ? current_field_num : field_num_8; // @[Serializerhw.scala 207:57 Serializerhw.scala 207:57 Serializerhw.scala 70:28]
  wire [5:0] _GEN_6214 = 4'h9 == stack_num ? current_field_num : field_num_9; // @[Serializerhw.scala 207:57 Serializerhw.scala 207:57 Serializerhw.scala 70:28]
  wire [5:0] _GEN_6215 = 4'ha == stack_num ? current_field_num : field_num_10; // @[Serializerhw.scala 207:57 Serializerhw.scala 207:57 Serializerhw.scala 70:28]
  wire [5:0] _GEN_6216 = 4'hb == stack_num ? current_field_num : field_num_11; // @[Serializerhw.scala 207:57 Serializerhw.scala 207:57 Serializerhw.scala 70:28]
  wire [5:0] _GEN_6217 = 4'hc == stack_num ? current_field_num : field_num_12; // @[Serializerhw.scala 207:57 Serializerhw.scala 207:57 Serializerhw.scala 70:28]
  wire [5:0] _GEN_6218 = 4'hd == stack_num ? current_field_num : field_num_13; // @[Serializerhw.scala 207:57 Serializerhw.scala 207:57 Serializerhw.scala 70:28]
  wire [5:0] _GEN_6219 = 4'he == stack_num ? current_field_num : field_num_14; // @[Serializerhw.scala 207:57 Serializerhw.scala 207:57 Serializerhw.scala 70:28]
  wire [5:0] _GEN_6220 = 4'hf == stack_num ? current_field_num : field_num_15; // @[Serializerhw.scala 207:57 Serializerhw.scala 207:57 Serializerhw.scala 70:28]
  wire [15:0] _GEN_6222 = c_sub_metadata_field_type == 5'hb ? c_sub_metadata_sub_class_id : 16'h0; // @[Serializerhw.scala 203:75 Serializerhw.scala 205:57 Util.scala 13:25]
  wire [3:0] _GEN_6223 = c_sub_metadata_field_type == 5'hb ? _stack_num_T_1 : stack_num; // @[Serializerhw.scala 203:75 Serializerhw.scala 206:57 Serializerhw.scala 76:30]
  wire [5:0] _GEN_6224 = c_sub_metadata_field_type == 5'hb ? _GEN_6205 : field_num_0; // @[Serializerhw.scala 203:75 Serializerhw.scala 70:28]
  wire [5:0] _GEN_6225 = c_sub_metadata_field_type == 5'hb ? _GEN_6206 : field_num_1; // @[Serializerhw.scala 203:75 Serializerhw.scala 70:28]
  wire [5:0] _GEN_6226 = c_sub_metadata_field_type == 5'hb ? _GEN_6207 : field_num_2; // @[Serializerhw.scala 203:75 Serializerhw.scala 70:28]
  wire [5:0] _GEN_6227 = c_sub_metadata_field_type == 5'hb ? _GEN_6208 : field_num_3; // @[Serializerhw.scala 203:75 Serializerhw.scala 70:28]
  wire [5:0] _GEN_6228 = c_sub_metadata_field_type == 5'hb ? _GEN_6209 : field_num_4; // @[Serializerhw.scala 203:75 Serializerhw.scala 70:28]
  wire [5:0] _GEN_6229 = c_sub_metadata_field_type == 5'hb ? _GEN_6210 : field_num_5; // @[Serializerhw.scala 203:75 Serializerhw.scala 70:28]
  wire [5:0] _GEN_6230 = c_sub_metadata_field_type == 5'hb ? _GEN_6211 : field_num_6; // @[Serializerhw.scala 203:75 Serializerhw.scala 70:28]
  wire [5:0] _GEN_6231 = c_sub_metadata_field_type == 5'hb ? _GEN_6212 : field_num_7; // @[Serializerhw.scala 203:75 Serializerhw.scala 70:28]
  wire [5:0] _GEN_6232 = c_sub_metadata_field_type == 5'hb ? _GEN_6213 : field_num_8; // @[Serializerhw.scala 203:75 Serializerhw.scala 70:28]
  wire [5:0] _GEN_6233 = c_sub_metadata_field_type == 5'hb ? _GEN_6214 : field_num_9; // @[Serializerhw.scala 203:75 Serializerhw.scala 70:28]
  wire [5:0] _GEN_6234 = c_sub_metadata_field_type == 5'hb ? _GEN_6215 : field_num_10; // @[Serializerhw.scala 203:75 Serializerhw.scala 70:28]
  wire [5:0] _GEN_6235 = c_sub_metadata_field_type == 5'hb ? _GEN_6216 : field_num_11; // @[Serializerhw.scala 203:75 Serializerhw.scala 70:28]
  wire [5:0] _GEN_6236 = c_sub_metadata_field_type == 5'hb ? _GEN_6217 : field_num_12; // @[Serializerhw.scala 203:75 Serializerhw.scala 70:28]
  wire [5:0] _GEN_6237 = c_sub_metadata_field_type == 5'hb ? _GEN_6218 : field_num_13; // @[Serializerhw.scala 203:75 Serializerhw.scala 70:28]
  wire [5:0] _GEN_6238 = c_sub_metadata_field_type == 5'hb ? _GEN_6219 : field_num_14; // @[Serializerhw.scala 203:75 Serializerhw.scala 70:28]
  wire [5:0] _GEN_6239 = c_sub_metadata_field_type == 5'hb ? _GEN_6220 : field_num_15; // @[Serializerhw.scala 203:75 Serializerhw.scala 70:28]
  wire [4:0] _GEN_6240 = c_sub_metadata_field_type == 5'hb ? 5'h11 : 5'hb; // @[Serializerhw.scala 203:75 Serializerhw.scala 208:57 Serializerhw.scala 211:53]
  wire [31:0] _GEN_6241 = c_sub_metadata_field_type == 5'hb ? current_field_length : {{16'd0},
    c_sub_metadata_sub_class_id}; // @[Serializerhw.scala 203:75 Serializerhw.scala 83:38 Serializerhw.scala 210:53]
  wire  _T_32 = 5'hb == state; // @[Conditional.scala 37:30]
  wire [31:0] _current_field_length_T_1 = current_field_length - 32'h1; // @[Serializerhw.scala 216:77]
  wire [31:0] _GEN_6242 = current_field_length > 32'h0 ? _current_field_length_T_1 : current_field_length; // @[Serializerhw.scala 215:43 Serializerhw.scala 216:53 Serializerhw.scala 83:38]
  wire [4:0] _GEN_6243 = current_field_length > 32'h0 ? 5'hb : 5'hc; // @[Serializerhw.scala 215:43 Serializerhw.scala 217:53 Serializerhw.scala 219:53]
  wire  _T_34 = 5'hc == state; // @[Conditional.scala 37:30]
  wire  _T_35 = 5'hd == state; // @[Conditional.scala 37:30]
  wire  _T_36 = 5'he == state; // @[Conditional.scala 37:30]
  wire [3:0] _current_field_num_T_11 = stack_num - 4'h1; // @[Serializerhw.scala 231:71]
  wire [5:0] _GEN_6261 = 4'h1 == _current_field_num_T_11 ? field_num_1 : field_num_0; // @[Serializerhw.scala 231:49 Serializerhw.scala 231:49]
  wire [5:0] _GEN_6262 = 4'h2 == _current_field_num_T_11 ? field_num_2 : _GEN_6261; // @[Serializerhw.scala 231:49 Serializerhw.scala 231:49]
  wire [5:0] _GEN_6263 = 4'h3 == _current_field_num_T_11 ? field_num_3 : _GEN_6262; // @[Serializerhw.scala 231:49 Serializerhw.scala 231:49]
  wire [5:0] _GEN_6264 = 4'h4 == _current_field_num_T_11 ? field_num_4 : _GEN_6263; // @[Serializerhw.scala 231:49 Serializerhw.scala 231:49]
  wire [5:0] _GEN_6265 = 4'h5 == _current_field_num_T_11 ? field_num_5 : _GEN_6264; // @[Serializerhw.scala 231:49 Serializerhw.scala 231:49]
  wire [5:0] _GEN_6266 = 4'h6 == _current_field_num_T_11 ? field_num_6 : _GEN_6265; // @[Serializerhw.scala 231:49 Serializerhw.scala 231:49]
  wire [5:0] _GEN_6267 = 4'h7 == _current_field_num_T_11 ? field_num_7 : _GEN_6266; // @[Serializerhw.scala 231:49 Serializerhw.scala 231:49]
  wire [5:0] _GEN_6268 = 4'h8 == _current_field_num_T_11 ? field_num_8 : _GEN_6267; // @[Serializerhw.scala 231:49 Serializerhw.scala 231:49]
  wire [5:0] _GEN_6269 = 4'h9 == _current_field_num_T_11 ? field_num_9 : _GEN_6268; // @[Serializerhw.scala 231:49 Serializerhw.scala 231:49]
  wire [5:0] _GEN_6270 = 4'ha == _current_field_num_T_11 ? field_num_10 : _GEN_6269; // @[Serializerhw.scala 231:49 Serializerhw.scala 231:49]
  wire [5:0] _GEN_6271 = 4'hb == _current_field_num_T_11 ? field_num_11 : _GEN_6270; // @[Serializerhw.scala 231:49 Serializerhw.scala 231:49]
  wire [5:0] _GEN_6272 = 4'hc == _current_field_num_T_11 ? field_num_12 : _GEN_6271; // @[Serializerhw.scala 231:49 Serializerhw.scala 231:49]
  wire [5:0] _GEN_6273 = 4'hd == _current_field_num_T_11 ? field_num_13 : _GEN_6272; // @[Serializerhw.scala 231:49 Serializerhw.scala 231:49]
  wire [5:0] _GEN_6274 = 4'he == _current_field_num_T_11 ? field_num_14 : _GEN_6273; // @[Serializerhw.scala 231:49 Serializerhw.scala 231:49]
  wire [5:0] _GEN_6275 = 4'hf == _current_field_num_T_11 ? field_num_15 : _GEN_6274; // @[Serializerhw.scala 231:49 Serializerhw.scala 231:49]
  wire  _T_37 = 5'hf == state; // @[Conditional.scala 37:30]
  wire  _T_38 = 5'h10 == state; // @[Conditional.scala 37:30]
  wire [4:0] _GEN_6278 = _T_38 ? 5'h6 : state; // @[Conditional.scala 39:67 Serializerhw.scala 242:49 Serializerhw.scala 86:46]
  wire [5:0] _GEN_6279 = _T_37 ? _current_field_num_T_1 : current_field_num; // @[Conditional.scala 39:67 Serializerhw.scala 236:49 Serializerhw.scala 73:36]
  wire [4:0] _GEN_6280 = _T_37 ? 5'h13 : _GEN_6278; // @[Conditional.scala 39:67 Serializerhw.scala 237:49]
  wire  _GEN_6281 = _T_37 ? 1'h0 : _T_38; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [5:0] _GEN_6283 = _T_36 ? _GEN_6205 : field_num_0; // @[Conditional.scala 39:67 Serializerhw.scala 70:28]
  wire [5:0] _GEN_6284 = _T_36 ? _GEN_6206 : field_num_1; // @[Conditional.scala 39:67 Serializerhw.scala 70:28]
  wire [5:0] _GEN_6285 = _T_36 ? _GEN_6207 : field_num_2; // @[Conditional.scala 39:67 Serializerhw.scala 70:28]
  wire [5:0] _GEN_6286 = _T_36 ? _GEN_6208 : field_num_3; // @[Conditional.scala 39:67 Serializerhw.scala 70:28]
  wire [5:0] _GEN_6287 = _T_36 ? _GEN_6209 : field_num_4; // @[Conditional.scala 39:67 Serializerhw.scala 70:28]
  wire [5:0] _GEN_6288 = _T_36 ? _GEN_6210 : field_num_5; // @[Conditional.scala 39:67 Serializerhw.scala 70:28]
  wire [5:0] _GEN_6289 = _T_36 ? _GEN_6211 : field_num_6; // @[Conditional.scala 39:67 Serializerhw.scala 70:28]
  wire [5:0] _GEN_6290 = _T_36 ? _GEN_6212 : field_num_7; // @[Conditional.scala 39:67 Serializerhw.scala 70:28]
  wire [5:0] _GEN_6291 = _T_36 ? _GEN_6213 : field_num_8; // @[Conditional.scala 39:67 Serializerhw.scala 70:28]
  wire [5:0] _GEN_6292 = _T_36 ? _GEN_6214 : field_num_9; // @[Conditional.scala 39:67 Serializerhw.scala 70:28]
  wire [5:0] _GEN_6293 = _T_36 ? _GEN_6215 : field_num_10; // @[Conditional.scala 39:67 Serializerhw.scala 70:28]
  wire [5:0] _GEN_6294 = _T_36 ? _GEN_6216 : field_num_11; // @[Conditional.scala 39:67 Serializerhw.scala 70:28]
  wire [5:0] _GEN_6295 = _T_36 ? _GEN_6217 : field_num_12; // @[Conditional.scala 39:67 Serializerhw.scala 70:28]
  wire [5:0] _GEN_6296 = _T_36 ? _GEN_6218 : field_num_13; // @[Conditional.scala 39:67 Serializerhw.scala 70:28]
  wire [5:0] _GEN_6297 = _T_36 ? _GEN_6219 : field_num_14; // @[Conditional.scala 39:67 Serializerhw.scala 70:28]
  wire [5:0] _GEN_6298 = _T_36 ? _GEN_6220 : field_num_15; // @[Conditional.scala 39:67 Serializerhw.scala 70:28]
  wire [5:0] _GEN_6299 = _T_36 ? _GEN_6275 : _GEN_6279; // @[Conditional.scala 39:67 Serializerhw.scala 231:49]
  wire [3:0] _GEN_6300 = _T_36 ? _current_field_num_T_11 : stack_num; // @[Conditional.scala 39:67 Serializerhw.scala 232:49 Serializerhw.scala 76:30]
  wire [4:0] _GEN_6301 = _T_36 ? 5'hd : _GEN_6280; // @[Conditional.scala 39:67 Serializerhw.scala 233:49]
  wire  _GEN_6302 = _T_36 ? 1'h0 : _GEN_6281; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [5:0] _GEN_6304 = _T_35 ? _current_field_num_T_1 : _GEN_6299; // @[Conditional.scala 39:67 Serializerhw.scala 226:49]
  wire [4:0] _GEN_6305 = _T_35 ? 5'h13 : _GEN_6301; // @[Conditional.scala 39:67 Serializerhw.scala 227:49]
  wire [5:0] _GEN_6306 = _T_35 ? field_num_0 : _GEN_6283; // @[Conditional.scala 39:67 Serializerhw.scala 70:28]
  wire [5:0] _GEN_6307 = _T_35 ? field_num_1 : _GEN_6284; // @[Conditional.scala 39:67 Serializerhw.scala 70:28]
  wire [5:0] _GEN_6308 = _T_35 ? field_num_2 : _GEN_6285; // @[Conditional.scala 39:67 Serializerhw.scala 70:28]
  wire [5:0] _GEN_6309 = _T_35 ? field_num_3 : _GEN_6286; // @[Conditional.scala 39:67 Serializerhw.scala 70:28]
  wire [5:0] _GEN_6310 = _T_35 ? field_num_4 : _GEN_6287; // @[Conditional.scala 39:67 Serializerhw.scala 70:28]
  wire [5:0] _GEN_6311 = _T_35 ? field_num_5 : _GEN_6288; // @[Conditional.scala 39:67 Serializerhw.scala 70:28]
  wire [5:0] _GEN_6312 = _T_35 ? field_num_6 : _GEN_6289; // @[Conditional.scala 39:67 Serializerhw.scala 70:28]
  wire [5:0] _GEN_6313 = _T_35 ? field_num_7 : _GEN_6290; // @[Conditional.scala 39:67 Serializerhw.scala 70:28]
  wire [5:0] _GEN_6314 = _T_35 ? field_num_8 : _GEN_6291; // @[Conditional.scala 39:67 Serializerhw.scala 70:28]
  wire [5:0] _GEN_6315 = _T_35 ? field_num_9 : _GEN_6292; // @[Conditional.scala 39:67 Serializerhw.scala 70:28]
  wire [5:0] _GEN_6316 = _T_35 ? field_num_10 : _GEN_6293; // @[Conditional.scala 39:67 Serializerhw.scala 70:28]
  wire [5:0] _GEN_6317 = _T_35 ? field_num_11 : _GEN_6294; // @[Conditional.scala 39:67 Serializerhw.scala 70:28]
  wire [5:0] _GEN_6318 = _T_35 ? field_num_12 : _GEN_6295; // @[Conditional.scala 39:67 Serializerhw.scala 70:28]
  wire [5:0] _GEN_6319 = _T_35 ? field_num_13 : _GEN_6296; // @[Conditional.scala 39:67 Serializerhw.scala 70:28]
  wire [5:0] _GEN_6320 = _T_35 ? field_num_14 : _GEN_6297; // @[Conditional.scala 39:67 Serializerhw.scala 70:28]
  wire [5:0] _GEN_6321 = _T_35 ? field_num_15 : _GEN_6298; // @[Conditional.scala 39:67 Serializerhw.scala 70:28]
  wire [3:0] _GEN_6322 = _T_35 ? stack_num : _GEN_6300; // @[Conditional.scala 39:67 Serializerhw.scala 76:30]
  wire  _GEN_6323 = _T_35 ? 1'h0 : _GEN_6302; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [4:0] _GEN_6325 = _T_34 ? 5'hd : _GEN_6305; // @[Conditional.scala 39:67 Serializerhw.scala 223:49]
  wire [5:0] _GEN_6326 = _T_34 ? current_field_num : _GEN_6304; // @[Conditional.scala 39:67 Serializerhw.scala 73:36]
  wire [5:0] _GEN_6327 = _T_34 ? field_num_0 : _GEN_6306; // @[Conditional.scala 39:67 Serializerhw.scala 70:28]
  wire [5:0] _GEN_6328 = _T_34 ? field_num_1 : _GEN_6307; // @[Conditional.scala 39:67 Serializerhw.scala 70:28]
  wire [5:0] _GEN_6329 = _T_34 ? field_num_2 : _GEN_6308; // @[Conditional.scala 39:67 Serializerhw.scala 70:28]
  wire [5:0] _GEN_6330 = _T_34 ? field_num_3 : _GEN_6309; // @[Conditional.scala 39:67 Serializerhw.scala 70:28]
  wire [5:0] _GEN_6331 = _T_34 ? field_num_4 : _GEN_6310; // @[Conditional.scala 39:67 Serializerhw.scala 70:28]
  wire [5:0] _GEN_6332 = _T_34 ? field_num_5 : _GEN_6311; // @[Conditional.scala 39:67 Serializerhw.scala 70:28]
  wire [5:0] _GEN_6333 = _T_34 ? field_num_6 : _GEN_6312; // @[Conditional.scala 39:67 Serializerhw.scala 70:28]
  wire [5:0] _GEN_6334 = _T_34 ? field_num_7 : _GEN_6313; // @[Conditional.scala 39:67 Serializerhw.scala 70:28]
  wire [5:0] _GEN_6335 = _T_34 ? field_num_8 : _GEN_6314; // @[Conditional.scala 39:67 Serializerhw.scala 70:28]
  wire [5:0] _GEN_6336 = _T_34 ? field_num_9 : _GEN_6315; // @[Conditional.scala 39:67 Serializerhw.scala 70:28]
  wire [5:0] _GEN_6337 = _T_34 ? field_num_10 : _GEN_6316; // @[Conditional.scala 39:67 Serializerhw.scala 70:28]
  wire [5:0] _GEN_6338 = _T_34 ? field_num_11 : _GEN_6317; // @[Conditional.scala 39:67 Serializerhw.scala 70:28]
  wire [5:0] _GEN_6339 = _T_34 ? field_num_12 : _GEN_6318; // @[Conditional.scala 39:67 Serializerhw.scala 70:28]
  wire [5:0] _GEN_6340 = _T_34 ? field_num_13 : _GEN_6319; // @[Conditional.scala 39:67 Serializerhw.scala 70:28]
  wire [5:0] _GEN_6341 = _T_34 ? field_num_14 : _GEN_6320; // @[Conditional.scala 39:67 Serializerhw.scala 70:28]
  wire [5:0] _GEN_6342 = _T_34 ? field_num_15 : _GEN_6321; // @[Conditional.scala 39:67 Serializerhw.scala 70:28]
  wire [3:0] _GEN_6343 = _T_34 ? stack_num : _GEN_6322; // @[Conditional.scala 39:67 Serializerhw.scala 76:30]
  wire  _GEN_6344 = _T_34 ? 1'h0 : _GEN_6323; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [31:0] _GEN_6346 = _T_32 ? _GEN_6242 : current_field_length; // @[Conditional.scala 39:67 Serializerhw.scala 83:38]
  wire [4:0] _GEN_6347 = _T_32 ? _GEN_6243 : _GEN_6325; // @[Conditional.scala 39:67]
  wire [5:0] _GEN_6348 = _T_32 ? current_field_num : _GEN_6326; // @[Conditional.scala 39:67 Serializerhw.scala 73:36]
  wire [5:0] _GEN_6349 = _T_32 ? field_num_0 : _GEN_6327; // @[Conditional.scala 39:67 Serializerhw.scala 70:28]
  wire [5:0] _GEN_6350 = _T_32 ? field_num_1 : _GEN_6328; // @[Conditional.scala 39:67 Serializerhw.scala 70:28]
  wire [5:0] _GEN_6351 = _T_32 ? field_num_2 : _GEN_6329; // @[Conditional.scala 39:67 Serializerhw.scala 70:28]
  wire [5:0] _GEN_6352 = _T_32 ? field_num_3 : _GEN_6330; // @[Conditional.scala 39:67 Serializerhw.scala 70:28]
  wire [5:0] _GEN_6353 = _T_32 ? field_num_4 : _GEN_6331; // @[Conditional.scala 39:67 Serializerhw.scala 70:28]
  wire [5:0] _GEN_6354 = _T_32 ? field_num_5 : _GEN_6332; // @[Conditional.scala 39:67 Serializerhw.scala 70:28]
  wire [5:0] _GEN_6355 = _T_32 ? field_num_6 : _GEN_6333; // @[Conditional.scala 39:67 Serializerhw.scala 70:28]
  wire [5:0] _GEN_6356 = _T_32 ? field_num_7 : _GEN_6334; // @[Conditional.scala 39:67 Serializerhw.scala 70:28]
  wire [5:0] _GEN_6357 = _T_32 ? field_num_8 : _GEN_6335; // @[Conditional.scala 39:67 Serializerhw.scala 70:28]
  wire [5:0] _GEN_6358 = _T_32 ? field_num_9 : _GEN_6336; // @[Conditional.scala 39:67 Serializerhw.scala 70:28]
  wire [5:0] _GEN_6359 = _T_32 ? field_num_10 : _GEN_6337; // @[Conditional.scala 39:67 Serializerhw.scala 70:28]
  wire [5:0] _GEN_6360 = _T_32 ? field_num_11 : _GEN_6338; // @[Conditional.scala 39:67 Serializerhw.scala 70:28]
  wire [5:0] _GEN_6361 = _T_32 ? field_num_12 : _GEN_6339; // @[Conditional.scala 39:67 Serializerhw.scala 70:28]
  wire [5:0] _GEN_6362 = _T_32 ? field_num_13 : _GEN_6340; // @[Conditional.scala 39:67 Serializerhw.scala 70:28]
  wire [5:0] _GEN_6363 = _T_32 ? field_num_14 : _GEN_6341; // @[Conditional.scala 39:67 Serializerhw.scala 70:28]
  wire [5:0] _GEN_6364 = _T_32 ? field_num_15 : _GEN_6342; // @[Conditional.scala 39:67 Serializerhw.scala 70:28]
  wire [3:0] _GEN_6365 = _T_32 ? stack_num : _GEN_6343; // @[Conditional.scala 39:67 Serializerhw.scala 76:30]
  wire  _GEN_6366 = _T_32 ? 1'h0 : _GEN_6344; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [15:0] _GEN_6369 = _T_30 ? _GEN_6222 : 16'h0; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [3:0] _GEN_6370 = _T_30 ? _GEN_6223 : _GEN_6365; // @[Conditional.scala 39:67]
  wire [5:0] _GEN_6371 = _T_30 ? _GEN_6224 : _GEN_6349; // @[Conditional.scala 39:67]
  wire [5:0] _GEN_6372 = _T_30 ? _GEN_6225 : _GEN_6350; // @[Conditional.scala 39:67]
  wire [5:0] _GEN_6373 = _T_30 ? _GEN_6226 : _GEN_6351; // @[Conditional.scala 39:67]
  wire [5:0] _GEN_6374 = _T_30 ? _GEN_6227 : _GEN_6352; // @[Conditional.scala 39:67]
  wire [5:0] _GEN_6375 = _T_30 ? _GEN_6228 : _GEN_6353; // @[Conditional.scala 39:67]
  wire [5:0] _GEN_6376 = _T_30 ? _GEN_6229 : _GEN_6354; // @[Conditional.scala 39:67]
  wire [5:0] _GEN_6377 = _T_30 ? _GEN_6230 : _GEN_6355; // @[Conditional.scala 39:67]
  wire [5:0] _GEN_6378 = _T_30 ? _GEN_6231 : _GEN_6356; // @[Conditional.scala 39:67]
  wire [5:0] _GEN_6379 = _T_30 ? _GEN_6232 : _GEN_6357; // @[Conditional.scala 39:67]
  wire [5:0] _GEN_6380 = _T_30 ? _GEN_6233 : _GEN_6358; // @[Conditional.scala 39:67]
  wire [5:0] _GEN_6381 = _T_30 ? _GEN_6234 : _GEN_6359; // @[Conditional.scala 39:67]
  wire [5:0] _GEN_6382 = _T_30 ? _GEN_6235 : _GEN_6360; // @[Conditional.scala 39:67]
  wire [5:0] _GEN_6383 = _T_30 ? _GEN_6236 : _GEN_6361; // @[Conditional.scala 39:67]
  wire [5:0] _GEN_6384 = _T_30 ? _GEN_6237 : _GEN_6362; // @[Conditional.scala 39:67]
  wire [5:0] _GEN_6385 = _T_30 ? _GEN_6238 : _GEN_6363; // @[Conditional.scala 39:67]
  wire [5:0] _GEN_6386 = _T_30 ? _GEN_6239 : _GEN_6364; // @[Conditional.scala 39:67]
  wire [4:0] _GEN_6387 = _T_30 ? _GEN_6240 : _GEN_6347; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_6388 = _T_30 ? _GEN_6241 : _GEN_6346; // @[Conditional.scala 39:67]
  wire [5:0] _GEN_6389 = _T_30 ? current_field_num : _GEN_6348; // @[Conditional.scala 39:67 Serializerhw.scala 73:36]
  wire  _GEN_6390 = _T_30 ? 1'h0 : _GEN_6366; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [4:0] _GEN_6392 = _T_27 ? _GEN_6202 : _GEN_6387; // @[Conditional.scala 39:67]
  wire [5:0] _GEN_6393 = _T_27 ? _GEN_6193 : _GEN_6389; // @[Conditional.scala 39:67]
  wire [7:0] _GEN_6394 = _T_27 ? _GEN_6194 : repeat_num; // @[Conditional.scala 39:67 Serializerhw.scala 75:29]
  wire  _GEN_6395 = _T_27 ? 1'h0 : _T_30 & _T_31; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [15:0] _GEN_6396 = _T_27 ? 16'h0 : _GEN_6369; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [3:0] _GEN_6397 = _T_27 ? stack_num : _GEN_6370; // @[Conditional.scala 39:67 Serializerhw.scala 76:30]
  wire [5:0] _GEN_6398 = _T_27 ? field_num_0 : _GEN_6371; // @[Conditional.scala 39:67 Serializerhw.scala 70:28]
  wire [5:0] _GEN_6399 = _T_27 ? field_num_1 : _GEN_6372; // @[Conditional.scala 39:67 Serializerhw.scala 70:28]
  wire [5:0] _GEN_6400 = _T_27 ? field_num_2 : _GEN_6373; // @[Conditional.scala 39:67 Serializerhw.scala 70:28]
  wire [5:0] _GEN_6401 = _T_27 ? field_num_3 : _GEN_6374; // @[Conditional.scala 39:67 Serializerhw.scala 70:28]
  wire [5:0] _GEN_6402 = _T_27 ? field_num_4 : _GEN_6375; // @[Conditional.scala 39:67 Serializerhw.scala 70:28]
  wire [5:0] _GEN_6403 = _T_27 ? field_num_5 : _GEN_6376; // @[Conditional.scala 39:67 Serializerhw.scala 70:28]
  wire [5:0] _GEN_6404 = _T_27 ? field_num_6 : _GEN_6377; // @[Conditional.scala 39:67 Serializerhw.scala 70:28]
  wire [5:0] _GEN_6405 = _T_27 ? field_num_7 : _GEN_6378; // @[Conditional.scala 39:67 Serializerhw.scala 70:28]
  wire [5:0] _GEN_6406 = _T_27 ? field_num_8 : _GEN_6379; // @[Conditional.scala 39:67 Serializerhw.scala 70:28]
  wire [5:0] _GEN_6407 = _T_27 ? field_num_9 : _GEN_6380; // @[Conditional.scala 39:67 Serializerhw.scala 70:28]
  wire [5:0] _GEN_6408 = _T_27 ? field_num_10 : _GEN_6381; // @[Conditional.scala 39:67 Serializerhw.scala 70:28]
  wire [5:0] _GEN_6409 = _T_27 ? field_num_11 : _GEN_6382; // @[Conditional.scala 39:67 Serializerhw.scala 70:28]
  wire [5:0] _GEN_6410 = _T_27 ? field_num_12 : _GEN_6383; // @[Conditional.scala 39:67 Serializerhw.scala 70:28]
  wire [5:0] _GEN_6411 = _T_27 ? field_num_13 : _GEN_6384; // @[Conditional.scala 39:67 Serializerhw.scala 70:28]
  wire [5:0] _GEN_6412 = _T_27 ? field_num_14 : _GEN_6385; // @[Conditional.scala 39:67 Serializerhw.scala 70:28]
  wire [5:0] _GEN_6413 = _T_27 ? field_num_15 : _GEN_6386; // @[Conditional.scala 39:67 Serializerhw.scala 70:28]
  wire [31:0] _GEN_6414 = _T_27 ? current_field_length : _GEN_6388; // @[Conditional.scala 39:67 Serializerhw.scala 83:38]
  wire  _GEN_6415 = _T_27 ? 1'h0 : _GEN_6390; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [4:0] _GEN_6417 = _T_24 ? _GEN_6197 : _GEN_6392; // @[Conditional.scala 39:67]
  wire [5:0] _GEN_6418 = _T_24 ? _GEN_6193 : _GEN_6393; // @[Conditional.scala 39:67]
  wire [7:0] _GEN_6419 = _T_24 ? _GEN_6194 : _GEN_6394; // @[Conditional.scala 39:67]
  wire  _GEN_6420 = _T_24 ? 1'h0 : _GEN_6395; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [15:0] _GEN_6421 = _T_24 ? 16'h0 : _GEN_6396; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [3:0] _GEN_6422 = _T_24 ? stack_num : _GEN_6397; // @[Conditional.scala 39:67 Serializerhw.scala 76:30]
  wire [5:0] _GEN_6423 = _T_24 ? field_num_0 : _GEN_6398; // @[Conditional.scala 39:67 Serializerhw.scala 70:28]
  wire [5:0] _GEN_6424 = _T_24 ? field_num_1 : _GEN_6399; // @[Conditional.scala 39:67 Serializerhw.scala 70:28]
  wire [5:0] _GEN_6425 = _T_24 ? field_num_2 : _GEN_6400; // @[Conditional.scala 39:67 Serializerhw.scala 70:28]
  wire [5:0] _GEN_6426 = _T_24 ? field_num_3 : _GEN_6401; // @[Conditional.scala 39:67 Serializerhw.scala 70:28]
  wire [5:0] _GEN_6427 = _T_24 ? field_num_4 : _GEN_6402; // @[Conditional.scala 39:67 Serializerhw.scala 70:28]
  wire [5:0] _GEN_6428 = _T_24 ? field_num_5 : _GEN_6403; // @[Conditional.scala 39:67 Serializerhw.scala 70:28]
  wire [5:0] _GEN_6429 = _T_24 ? field_num_6 : _GEN_6404; // @[Conditional.scala 39:67 Serializerhw.scala 70:28]
  wire [5:0] _GEN_6430 = _T_24 ? field_num_7 : _GEN_6405; // @[Conditional.scala 39:67 Serializerhw.scala 70:28]
  wire [5:0] _GEN_6431 = _T_24 ? field_num_8 : _GEN_6406; // @[Conditional.scala 39:67 Serializerhw.scala 70:28]
  wire [5:0] _GEN_6432 = _T_24 ? field_num_9 : _GEN_6407; // @[Conditional.scala 39:67 Serializerhw.scala 70:28]
  wire [5:0] _GEN_6433 = _T_24 ? field_num_10 : _GEN_6408; // @[Conditional.scala 39:67 Serializerhw.scala 70:28]
  wire [5:0] _GEN_6434 = _T_24 ? field_num_11 : _GEN_6409; // @[Conditional.scala 39:67 Serializerhw.scala 70:28]
  wire [5:0] _GEN_6435 = _T_24 ? field_num_12 : _GEN_6410; // @[Conditional.scala 39:67 Serializerhw.scala 70:28]
  wire [5:0] _GEN_6436 = _T_24 ? field_num_13 : _GEN_6411; // @[Conditional.scala 39:67 Serializerhw.scala 70:28]
  wire [5:0] _GEN_6437 = _T_24 ? field_num_14 : _GEN_6412; // @[Conditional.scala 39:67 Serializerhw.scala 70:28]
  wire [5:0] _GEN_6438 = _T_24 ? field_num_15 : _GEN_6413; // @[Conditional.scala 39:67 Serializerhw.scala 70:28]
  wire [31:0] _GEN_6439 = _T_24 ? current_field_length : _GEN_6414; // @[Conditional.scala 39:67 Serializerhw.scala 83:38]
  wire  _GEN_6440 = _T_24 ? 1'h0 : _GEN_6415; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [4:0] _GEN_6442 = _T_21 ? _GEN_6192 : _GEN_6417; // @[Conditional.scala 39:67]
  wire [5:0] _GEN_6443 = _T_21 ? _GEN_6193 : _GEN_6418; // @[Conditional.scala 39:67]
  wire [7:0] _GEN_6444 = _T_21 ? _GEN_6194 : _GEN_6419; // @[Conditional.scala 39:67]
  wire  _GEN_6445 = _T_21 ? 1'h0 : _GEN_6420; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [15:0] _GEN_6446 = _T_21 ? 16'h0 : _GEN_6421; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [3:0] _GEN_6447 = _T_21 ? stack_num : _GEN_6422; // @[Conditional.scala 39:67 Serializerhw.scala 76:30]
  wire [5:0] _GEN_6448 = _T_21 ? field_num_0 : _GEN_6423; // @[Conditional.scala 39:67 Serializerhw.scala 70:28]
  wire [5:0] _GEN_6449 = _T_21 ? field_num_1 : _GEN_6424; // @[Conditional.scala 39:67 Serializerhw.scala 70:28]
  wire [5:0] _GEN_6450 = _T_21 ? field_num_2 : _GEN_6425; // @[Conditional.scala 39:67 Serializerhw.scala 70:28]
  wire [5:0] _GEN_6451 = _T_21 ? field_num_3 : _GEN_6426; // @[Conditional.scala 39:67 Serializerhw.scala 70:28]
  wire [5:0] _GEN_6452 = _T_21 ? field_num_4 : _GEN_6427; // @[Conditional.scala 39:67 Serializerhw.scala 70:28]
  wire [5:0] _GEN_6453 = _T_21 ? field_num_5 : _GEN_6428; // @[Conditional.scala 39:67 Serializerhw.scala 70:28]
  wire [5:0] _GEN_6454 = _T_21 ? field_num_6 : _GEN_6429; // @[Conditional.scala 39:67 Serializerhw.scala 70:28]
  wire [5:0] _GEN_6455 = _T_21 ? field_num_7 : _GEN_6430; // @[Conditional.scala 39:67 Serializerhw.scala 70:28]
  wire [5:0] _GEN_6456 = _T_21 ? field_num_8 : _GEN_6431; // @[Conditional.scala 39:67 Serializerhw.scala 70:28]
  wire [5:0] _GEN_6457 = _T_21 ? field_num_9 : _GEN_6432; // @[Conditional.scala 39:67 Serializerhw.scala 70:28]
  wire [5:0] _GEN_6458 = _T_21 ? field_num_10 : _GEN_6433; // @[Conditional.scala 39:67 Serializerhw.scala 70:28]
  wire [5:0] _GEN_6459 = _T_21 ? field_num_11 : _GEN_6434; // @[Conditional.scala 39:67 Serializerhw.scala 70:28]
  wire [5:0] _GEN_6460 = _T_21 ? field_num_12 : _GEN_6435; // @[Conditional.scala 39:67 Serializerhw.scala 70:28]
  wire [5:0] _GEN_6461 = _T_21 ? field_num_13 : _GEN_6436; // @[Conditional.scala 39:67 Serializerhw.scala 70:28]
  wire [5:0] _GEN_6462 = _T_21 ? field_num_14 : _GEN_6437; // @[Conditional.scala 39:67 Serializerhw.scala 70:28]
  wire [5:0] _GEN_6463 = _T_21 ? field_num_15 : _GEN_6438; // @[Conditional.scala 39:67 Serializerhw.scala 70:28]
  wire [31:0] _GEN_6464 = _T_21 ? current_field_length : _GEN_6439; // @[Conditional.scala 39:67 Serializerhw.scala 83:38]
  wire  _GEN_6465 = _T_21 ? 1'h0 : _GEN_6440; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [15:0] _GEN_6467 = _T_14 ? _GEN_6188 : {{8'd0}, _GEN_6444}; // @[Conditional.scala 39:67]
  wire [4:0] _GEN_6468 = _T_14 ? _GEN_6189 : _GEN_6442; // @[Conditional.scala 39:67]
  wire [5:0] _GEN_6469 = _T_14 ? current_field_num : _GEN_6443; // @[Conditional.scala 39:67 Serializerhw.scala 73:36]
  wire  _GEN_6470 = _T_14 ? 1'h0 : _GEN_6445; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [15:0] _GEN_6471 = _T_14 ? 16'h0 : _GEN_6446; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [3:0] _GEN_6472 = _T_14 ? stack_num : _GEN_6447; // @[Conditional.scala 39:67 Serializerhw.scala 76:30]
  wire [5:0] _GEN_6473 = _T_14 ? field_num_0 : _GEN_6448; // @[Conditional.scala 39:67 Serializerhw.scala 70:28]
  wire [5:0] _GEN_6474 = _T_14 ? field_num_1 : _GEN_6449; // @[Conditional.scala 39:67 Serializerhw.scala 70:28]
  wire [5:0] _GEN_6475 = _T_14 ? field_num_2 : _GEN_6450; // @[Conditional.scala 39:67 Serializerhw.scala 70:28]
  wire [5:0] _GEN_6476 = _T_14 ? field_num_3 : _GEN_6451; // @[Conditional.scala 39:67 Serializerhw.scala 70:28]
  wire [5:0] _GEN_6477 = _T_14 ? field_num_4 : _GEN_6452; // @[Conditional.scala 39:67 Serializerhw.scala 70:28]
  wire [5:0] _GEN_6478 = _T_14 ? field_num_5 : _GEN_6453; // @[Conditional.scala 39:67 Serializerhw.scala 70:28]
  wire [5:0] _GEN_6479 = _T_14 ? field_num_6 : _GEN_6454; // @[Conditional.scala 39:67 Serializerhw.scala 70:28]
  wire [5:0] _GEN_6480 = _T_14 ? field_num_7 : _GEN_6455; // @[Conditional.scala 39:67 Serializerhw.scala 70:28]
  wire [5:0] _GEN_6481 = _T_14 ? field_num_8 : _GEN_6456; // @[Conditional.scala 39:67 Serializerhw.scala 70:28]
  wire [5:0] _GEN_6482 = _T_14 ? field_num_9 : _GEN_6457; // @[Conditional.scala 39:67 Serializerhw.scala 70:28]
  wire [5:0] _GEN_6483 = _T_14 ? field_num_10 : _GEN_6458; // @[Conditional.scala 39:67 Serializerhw.scala 70:28]
  wire [5:0] _GEN_6484 = _T_14 ? field_num_11 : _GEN_6459; // @[Conditional.scala 39:67 Serializerhw.scala 70:28]
  wire [5:0] _GEN_6485 = _T_14 ? field_num_12 : _GEN_6460; // @[Conditional.scala 39:67 Serializerhw.scala 70:28]
  wire [5:0] _GEN_6486 = _T_14 ? field_num_13 : _GEN_6461; // @[Conditional.scala 39:67 Serializerhw.scala 70:28]
  wire [5:0] _GEN_6487 = _T_14 ? field_num_14 : _GEN_6462; // @[Conditional.scala 39:67 Serializerhw.scala 70:28]
  wire [5:0] _GEN_6488 = _T_14 ? field_num_15 : _GEN_6463; // @[Conditional.scala 39:67 Serializerhw.scala 70:28]
  wire [31:0] _GEN_6489 = _T_14 ? current_field_length : _GEN_6464; // @[Conditional.scala 39:67 Serializerhw.scala 83:38]
  wire  _GEN_6490 = _T_14 ? 1'h0 : _GEN_6465; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [4:0] _GEN_6492 = _T_10 ? _GEN_6062 : _GEN_6468; // @[Conditional.scala 39:67]
  wire [5:0] _GEN_6493 = _T_10 ? _GEN_6063 : _GEN_6469; // @[Conditional.scala 39:67]
  wire [15:0] _GEN_6495 = _T_10 ? _GEN_6065 : c_sub_metadata_sub_class_id; // @[Conditional.scala 39:67 Serializerhw.scala 74:33]
  wire [4:0] _GEN_6496 = _T_10 ? _GEN_6066 : c_sub_metadata_field_type; // @[Conditional.scala 39:67 Serializerhw.scala 74:33]
  wire  _GEN_6497 = _T_10 ? _GEN_6067 : c_sub_metadata_is_repeated; // @[Conditional.scala 39:67 Serializerhw.scala 74:33]
  wire [15:0] _GEN_6498 = _T_10 ? {{8'd0}, repeat_num} : _GEN_6467; // @[Conditional.scala 39:67 Serializerhw.scala 75:29]
  wire  _GEN_6499 = _T_10 ? 1'h0 : _GEN_6470; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [15:0] _GEN_6500 = _T_10 ? 16'h0 : _GEN_6471; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [3:0] _GEN_6501 = _T_10 ? stack_num : _GEN_6472; // @[Conditional.scala 39:67 Serializerhw.scala 76:30]
  wire [5:0] _GEN_6502 = _T_10 ? field_num_0 : _GEN_6473; // @[Conditional.scala 39:67 Serializerhw.scala 70:28]
  wire [5:0] _GEN_6503 = _T_10 ? field_num_1 : _GEN_6474; // @[Conditional.scala 39:67 Serializerhw.scala 70:28]
  wire [5:0] _GEN_6504 = _T_10 ? field_num_2 : _GEN_6475; // @[Conditional.scala 39:67 Serializerhw.scala 70:28]
  wire [5:0] _GEN_6505 = _T_10 ? field_num_3 : _GEN_6476; // @[Conditional.scala 39:67 Serializerhw.scala 70:28]
  wire [5:0] _GEN_6506 = _T_10 ? field_num_4 : _GEN_6477; // @[Conditional.scala 39:67 Serializerhw.scala 70:28]
  wire [5:0] _GEN_6507 = _T_10 ? field_num_5 : _GEN_6478; // @[Conditional.scala 39:67 Serializerhw.scala 70:28]
  wire [5:0] _GEN_6508 = _T_10 ? field_num_6 : _GEN_6479; // @[Conditional.scala 39:67 Serializerhw.scala 70:28]
  wire [5:0] _GEN_6509 = _T_10 ? field_num_7 : _GEN_6480; // @[Conditional.scala 39:67 Serializerhw.scala 70:28]
  wire [5:0] _GEN_6510 = _T_10 ? field_num_8 : _GEN_6481; // @[Conditional.scala 39:67 Serializerhw.scala 70:28]
  wire [5:0] _GEN_6511 = _T_10 ? field_num_9 : _GEN_6482; // @[Conditional.scala 39:67 Serializerhw.scala 70:28]
  wire [5:0] _GEN_6512 = _T_10 ? field_num_10 : _GEN_6483; // @[Conditional.scala 39:67 Serializerhw.scala 70:28]
  wire [5:0] _GEN_6513 = _T_10 ? field_num_11 : _GEN_6484; // @[Conditional.scala 39:67 Serializerhw.scala 70:28]
  wire [5:0] _GEN_6514 = _T_10 ? field_num_12 : _GEN_6485; // @[Conditional.scala 39:67 Serializerhw.scala 70:28]
  wire [5:0] _GEN_6515 = _T_10 ? field_num_13 : _GEN_6486; // @[Conditional.scala 39:67 Serializerhw.scala 70:28]
  wire [5:0] _GEN_6516 = _T_10 ? field_num_14 : _GEN_6487; // @[Conditional.scala 39:67 Serializerhw.scala 70:28]
  wire [5:0] _GEN_6517 = _T_10 ? field_num_15 : _GEN_6488; // @[Conditional.scala 39:67 Serializerhw.scala 70:28]
  wire [31:0] _GEN_6518 = _T_10 ? current_field_length : _GEN_6489; // @[Conditional.scala 39:67 Serializerhw.scala 83:38]
  wire  _GEN_6519 = _T_10 ? 1'h0 : _GEN_6490; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [5:0] _GEN_6522 = _T_8 ? current_field_num : _GEN_6493; // @[Conditional.scala 39:67 Serializerhw.scala 73:36]
  wire [15:0] _GEN_6527 = _T_8 ? {{8'd0}, repeat_num} : _GEN_6498; // @[Conditional.scala 39:67 Serializerhw.scala 75:29]
  wire  _GEN_6528 = _T_8 ? 1'h0 : _GEN_6499; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [15:0] _GEN_6529 = _T_8 ? 16'h0 : _GEN_6500; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire  _GEN_6548 = _T_8 ? 1'h0 : _GEN_6519; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [7:0] _GEN_8576 = _T_6 ? _GEN_4068 : {{2'd0}, _GEN_6522}; // @[Conditional.scala 39:67]
  wire  _GEN_8578 = _T_6 & _T_7; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [63:0] _GEN_8579 = _T_6 ? _GEN_4071 : 64'h0; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [31:0] _GEN_8580 = _T_6 ? _GEN_4072 : 32'h0; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [15:0] _GEN_8586 = _T_6 ? {{8'd0}, repeat_num} : _GEN_6527; // @[Conditional.scala 39:67 Serializerhw.scala 75:29]
  wire  _GEN_8587 = _T_6 ? 1'h0 : _GEN_6528; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [15:0] _GEN_8588 = _T_6 ? 16'h0 : _GEN_6529; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire  _GEN_8591 = _T_6 ? 1'h0 : _GEN_6548; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [15:0] _GEN_8601 = _T_4 ? {{6'd0}, _GEN_12} : _GEN_8588; // @[Conditional.scala 40:58]
  wire [7:0] _GEN_10631 = _T_4 ? {{2'd0}, current_field_num} : _GEN_8576; // @[Conditional.scala 40:58 Serializerhw.scala 73:36]
  wire [15:0] _GEN_10639 = _T_4 ? {{8'd0}, repeat_num} : _GEN_8586; // @[Conditional.scala 40:58 Serializerhw.scala 75:29]
  XQueue_2 meta_in_fifo ( // @[XQueue.scala 35:23]
    .clock(meta_in_fifo_clock),
    .reset(meta_in_fifo_reset),
    .io_in_ready(meta_in_fifo_io_in_ready),
    .io_in_valid(meta_in_fifo_io_in_valid),
    .io_in_bits_class_id(meta_in_fifo_io_in_bits_class_id),
    .io_in_bits_host_base_addr(meta_in_fifo_io_in_bits_host_base_addr),
    .io_out_ready(meta_in_fifo_io_out_ready),
    .io_out_valid(meta_in_fifo_io_out_valid),
    .io_out_bits_class_id(meta_in_fifo_io_out_bits_class_id),
    .io_out_bits_host_base_addr(meta_in_fifo_io_out_bits_host_base_addr)
  );
  XQueue_3 class_meta_rsp_fifo ( // @[XQueue.scala 35:23]
    .clock(class_meta_rsp_fifo_clock),
    .reset(class_meta_rsp_fifo_reset),
    .io_in_valid(class_meta_rsp_fifo_io_in_valid),
    .io_in_bits_class_meta_max_field_num(class_meta_rsp_fifo_io_in_bits_class_meta_max_field_num),
    .io_in_bits_class_meta_field_type_0_is_repeated(class_meta_rsp_fifo_io_in_bits_class_meta_field_type_0_is_repeated),
    .io_in_bits_class_meta_field_type_0_field_type(class_meta_rsp_fifo_io_in_bits_class_meta_field_type_0_field_type),
    .io_in_bits_class_meta_field_type_0_sub_class_id(class_meta_rsp_fifo_io_in_bits_class_meta_field_type_0_sub_class_id
      ),
    .io_in_bits_class_meta_field_type_1_is_repeated(class_meta_rsp_fifo_io_in_bits_class_meta_field_type_1_is_repeated),
    .io_in_bits_class_meta_field_type_1_field_type(class_meta_rsp_fifo_io_in_bits_class_meta_field_type_1_field_type),
    .io_in_bits_class_meta_field_type_1_sub_class_id(class_meta_rsp_fifo_io_in_bits_class_meta_field_type_1_sub_class_id
      ),
    .io_in_bits_class_meta_field_type_2_is_repeated(class_meta_rsp_fifo_io_in_bits_class_meta_field_type_2_is_repeated),
    .io_in_bits_class_meta_field_type_2_field_type(class_meta_rsp_fifo_io_in_bits_class_meta_field_type_2_field_type),
    .io_in_bits_class_meta_field_type_2_sub_class_id(class_meta_rsp_fifo_io_in_bits_class_meta_field_type_2_sub_class_id
      ),
    .io_in_bits_class_meta_field_type_3_is_repeated(class_meta_rsp_fifo_io_in_bits_class_meta_field_type_3_is_repeated),
    .io_in_bits_class_meta_field_type_3_field_type(class_meta_rsp_fifo_io_in_bits_class_meta_field_type_3_field_type),
    .io_in_bits_class_meta_field_type_3_sub_class_id(class_meta_rsp_fifo_io_in_bits_class_meta_field_type_3_sub_class_id
      ),
    .io_in_bits_class_meta_field_type_4_is_repeated(class_meta_rsp_fifo_io_in_bits_class_meta_field_type_4_is_repeated),
    .io_in_bits_class_meta_field_type_4_field_type(class_meta_rsp_fifo_io_in_bits_class_meta_field_type_4_field_type),
    .io_in_bits_class_meta_field_type_4_sub_class_id(class_meta_rsp_fifo_io_in_bits_class_meta_field_type_4_sub_class_id
      ),
    .io_in_bits_class_meta_field_type_5_is_repeated(class_meta_rsp_fifo_io_in_bits_class_meta_field_type_5_is_repeated),
    .io_in_bits_class_meta_field_type_5_field_type(class_meta_rsp_fifo_io_in_bits_class_meta_field_type_5_field_type),
    .io_in_bits_class_meta_field_type_5_sub_class_id(class_meta_rsp_fifo_io_in_bits_class_meta_field_type_5_sub_class_id
      ),
    .io_in_bits_class_meta_field_type_6_is_repeated(class_meta_rsp_fifo_io_in_bits_class_meta_field_type_6_is_repeated),
    .io_in_bits_class_meta_field_type_6_field_type(class_meta_rsp_fifo_io_in_bits_class_meta_field_type_6_field_type),
    .io_in_bits_class_meta_field_type_6_sub_class_id(class_meta_rsp_fifo_io_in_bits_class_meta_field_type_6_sub_class_id
      ),
    .io_in_bits_class_meta_field_type_7_is_repeated(class_meta_rsp_fifo_io_in_bits_class_meta_field_type_7_is_repeated),
    .io_in_bits_class_meta_field_type_7_field_type(class_meta_rsp_fifo_io_in_bits_class_meta_field_type_7_field_type),
    .io_in_bits_class_meta_field_type_7_sub_class_id(class_meta_rsp_fifo_io_in_bits_class_meta_field_type_7_sub_class_id
      ),
    .io_in_bits_class_meta_field_type_8_is_repeated(class_meta_rsp_fifo_io_in_bits_class_meta_field_type_8_is_repeated),
    .io_in_bits_class_meta_field_type_8_field_type(class_meta_rsp_fifo_io_in_bits_class_meta_field_type_8_field_type),
    .io_in_bits_class_meta_field_type_8_sub_class_id(class_meta_rsp_fifo_io_in_bits_class_meta_field_type_8_sub_class_id
      ),
    .io_in_bits_class_meta_field_type_9_is_repeated(class_meta_rsp_fifo_io_in_bits_class_meta_field_type_9_is_repeated),
    .io_in_bits_class_meta_field_type_9_field_type(class_meta_rsp_fifo_io_in_bits_class_meta_field_type_9_field_type),
    .io_in_bits_class_meta_field_type_9_sub_class_id(class_meta_rsp_fifo_io_in_bits_class_meta_field_type_9_sub_class_id
      ),
    .io_in_bits_class_meta_field_type_10_is_repeated(class_meta_rsp_fifo_io_in_bits_class_meta_field_type_10_is_repeated
      ),
    .io_in_bits_class_meta_field_type_10_field_type(class_meta_rsp_fifo_io_in_bits_class_meta_field_type_10_field_type),
    .io_in_bits_class_meta_field_type_10_sub_class_id(
      class_meta_rsp_fifo_io_in_bits_class_meta_field_type_10_sub_class_id),
    .io_in_bits_class_meta_field_type_11_is_repeated(class_meta_rsp_fifo_io_in_bits_class_meta_field_type_11_is_repeated
      ),
    .io_in_bits_class_meta_field_type_11_field_type(class_meta_rsp_fifo_io_in_bits_class_meta_field_type_11_field_type),
    .io_in_bits_class_meta_field_type_11_sub_class_id(
      class_meta_rsp_fifo_io_in_bits_class_meta_field_type_11_sub_class_id),
    .io_in_bits_class_meta_field_type_12_is_repeated(class_meta_rsp_fifo_io_in_bits_class_meta_field_type_12_is_repeated
      ),
    .io_in_bits_class_meta_field_type_12_field_type(class_meta_rsp_fifo_io_in_bits_class_meta_field_type_12_field_type),
    .io_in_bits_class_meta_field_type_12_sub_class_id(
      class_meta_rsp_fifo_io_in_bits_class_meta_field_type_12_sub_class_id),
    .io_in_bits_class_meta_field_type_13_is_repeated(class_meta_rsp_fifo_io_in_bits_class_meta_field_type_13_is_repeated
      ),
    .io_in_bits_class_meta_field_type_13_field_type(class_meta_rsp_fifo_io_in_bits_class_meta_field_type_13_field_type),
    .io_in_bits_class_meta_field_type_13_sub_class_id(
      class_meta_rsp_fifo_io_in_bits_class_meta_field_type_13_sub_class_id),
    .io_in_bits_class_meta_field_type_14_is_repeated(class_meta_rsp_fifo_io_in_bits_class_meta_field_type_14_is_repeated
      ),
    .io_in_bits_class_meta_field_type_14_field_type(class_meta_rsp_fifo_io_in_bits_class_meta_field_type_14_field_type),
    .io_in_bits_class_meta_field_type_14_sub_class_id(
      class_meta_rsp_fifo_io_in_bits_class_meta_field_type_14_sub_class_id),
    .io_in_bits_class_meta_field_type_15_is_repeated(class_meta_rsp_fifo_io_in_bits_class_meta_field_type_15_is_repeated
      ),
    .io_in_bits_class_meta_field_type_15_field_type(class_meta_rsp_fifo_io_in_bits_class_meta_field_type_15_field_type),
    .io_in_bits_class_meta_field_type_15_sub_class_id(
      class_meta_rsp_fifo_io_in_bits_class_meta_field_type_15_sub_class_id),
    .io_in_bits_class_meta_field_type_16_is_repeated(class_meta_rsp_fifo_io_in_bits_class_meta_field_type_16_is_repeated
      ),
    .io_in_bits_class_meta_field_type_16_field_type(class_meta_rsp_fifo_io_in_bits_class_meta_field_type_16_field_type),
    .io_in_bits_class_meta_field_type_16_sub_class_id(
      class_meta_rsp_fifo_io_in_bits_class_meta_field_type_16_sub_class_id),
    .io_in_bits_class_meta_field_type_17_is_repeated(class_meta_rsp_fifo_io_in_bits_class_meta_field_type_17_is_repeated
      ),
    .io_in_bits_class_meta_field_type_17_field_type(class_meta_rsp_fifo_io_in_bits_class_meta_field_type_17_field_type),
    .io_in_bits_class_meta_field_type_17_sub_class_id(
      class_meta_rsp_fifo_io_in_bits_class_meta_field_type_17_sub_class_id),
    .io_in_bits_class_meta_field_type_18_is_repeated(class_meta_rsp_fifo_io_in_bits_class_meta_field_type_18_is_repeated
      ),
    .io_in_bits_class_meta_field_type_18_field_type(class_meta_rsp_fifo_io_in_bits_class_meta_field_type_18_field_type),
    .io_in_bits_class_meta_field_type_18_sub_class_id(
      class_meta_rsp_fifo_io_in_bits_class_meta_field_type_18_sub_class_id),
    .io_in_bits_class_meta_field_type_19_is_repeated(class_meta_rsp_fifo_io_in_bits_class_meta_field_type_19_is_repeated
      ),
    .io_in_bits_class_meta_field_type_19_field_type(class_meta_rsp_fifo_io_in_bits_class_meta_field_type_19_field_type),
    .io_in_bits_class_meta_field_type_19_sub_class_id(
      class_meta_rsp_fifo_io_in_bits_class_meta_field_type_19_sub_class_id),
    .io_in_bits_class_meta_field_type_20_is_repeated(class_meta_rsp_fifo_io_in_bits_class_meta_field_type_20_is_repeated
      ),
    .io_in_bits_class_meta_field_type_20_field_type(class_meta_rsp_fifo_io_in_bits_class_meta_field_type_20_field_type),
    .io_in_bits_class_meta_field_type_20_sub_class_id(
      class_meta_rsp_fifo_io_in_bits_class_meta_field_type_20_sub_class_id),
    .io_in_bits_class_meta_field_type_21_is_repeated(class_meta_rsp_fifo_io_in_bits_class_meta_field_type_21_is_repeated
      ),
    .io_in_bits_class_meta_field_type_21_field_type(class_meta_rsp_fifo_io_in_bits_class_meta_field_type_21_field_type),
    .io_in_bits_class_meta_field_type_21_sub_class_id(
      class_meta_rsp_fifo_io_in_bits_class_meta_field_type_21_sub_class_id),
    .io_in_bits_class_meta_field_type_22_is_repeated(class_meta_rsp_fifo_io_in_bits_class_meta_field_type_22_is_repeated
      ),
    .io_in_bits_class_meta_field_type_22_field_type(class_meta_rsp_fifo_io_in_bits_class_meta_field_type_22_field_type),
    .io_in_bits_class_meta_field_type_22_sub_class_id(
      class_meta_rsp_fifo_io_in_bits_class_meta_field_type_22_sub_class_id),
    .io_in_bits_class_meta_field_type_23_is_repeated(class_meta_rsp_fifo_io_in_bits_class_meta_field_type_23_is_repeated
      ),
    .io_in_bits_class_meta_field_type_23_field_type(class_meta_rsp_fifo_io_in_bits_class_meta_field_type_23_field_type),
    .io_in_bits_class_meta_field_type_23_sub_class_id(
      class_meta_rsp_fifo_io_in_bits_class_meta_field_type_23_sub_class_id),
    .io_in_bits_class_meta_field_type_24_is_repeated(class_meta_rsp_fifo_io_in_bits_class_meta_field_type_24_is_repeated
      ),
    .io_in_bits_class_meta_field_type_24_field_type(class_meta_rsp_fifo_io_in_bits_class_meta_field_type_24_field_type),
    .io_in_bits_class_meta_field_type_24_sub_class_id(
      class_meta_rsp_fifo_io_in_bits_class_meta_field_type_24_sub_class_id),
    .io_in_bits_class_meta_field_type_25_is_repeated(class_meta_rsp_fifo_io_in_bits_class_meta_field_type_25_is_repeated
      ),
    .io_in_bits_class_meta_field_type_25_field_type(class_meta_rsp_fifo_io_in_bits_class_meta_field_type_25_field_type),
    .io_in_bits_class_meta_field_type_25_sub_class_id(
      class_meta_rsp_fifo_io_in_bits_class_meta_field_type_25_sub_class_id),
    .io_in_bits_class_meta_field_type_26_is_repeated(class_meta_rsp_fifo_io_in_bits_class_meta_field_type_26_is_repeated
      ),
    .io_in_bits_class_meta_field_type_26_field_type(class_meta_rsp_fifo_io_in_bits_class_meta_field_type_26_field_type),
    .io_in_bits_class_meta_field_type_26_sub_class_id(
      class_meta_rsp_fifo_io_in_bits_class_meta_field_type_26_sub_class_id),
    .io_in_bits_class_meta_field_type_27_is_repeated(class_meta_rsp_fifo_io_in_bits_class_meta_field_type_27_is_repeated
      ),
    .io_in_bits_class_meta_field_type_27_field_type(class_meta_rsp_fifo_io_in_bits_class_meta_field_type_27_field_type),
    .io_in_bits_class_meta_field_type_27_sub_class_id(
      class_meta_rsp_fifo_io_in_bits_class_meta_field_type_27_sub_class_id),
    .io_in_bits_class_meta_field_type_28_is_repeated(class_meta_rsp_fifo_io_in_bits_class_meta_field_type_28_is_repeated
      ),
    .io_in_bits_class_meta_field_type_28_field_type(class_meta_rsp_fifo_io_in_bits_class_meta_field_type_28_field_type),
    .io_in_bits_class_meta_field_type_28_sub_class_id(
      class_meta_rsp_fifo_io_in_bits_class_meta_field_type_28_sub_class_id),
    .io_in_bits_class_meta_field_type_29_is_repeated(class_meta_rsp_fifo_io_in_bits_class_meta_field_type_29_is_repeated
      ),
    .io_in_bits_class_meta_field_type_29_field_type(class_meta_rsp_fifo_io_in_bits_class_meta_field_type_29_field_type),
    .io_in_bits_class_meta_field_type_29_sub_class_id(
      class_meta_rsp_fifo_io_in_bits_class_meta_field_type_29_sub_class_id),
    .io_in_bits_class_meta_field_type_30_is_repeated(class_meta_rsp_fifo_io_in_bits_class_meta_field_type_30_is_repeated
      ),
    .io_in_bits_class_meta_field_type_30_field_type(class_meta_rsp_fifo_io_in_bits_class_meta_field_type_30_field_type),
    .io_in_bits_class_meta_field_type_30_sub_class_id(
      class_meta_rsp_fifo_io_in_bits_class_meta_field_type_30_sub_class_id),
    .io_in_bits_class_meta_field_type_31_is_repeated(class_meta_rsp_fifo_io_in_bits_class_meta_field_type_31_is_repeated
      ),
    .io_in_bits_class_meta_field_type_31_field_type(class_meta_rsp_fifo_io_in_bits_class_meta_field_type_31_field_type),
    .io_in_bits_class_meta_field_type_31_sub_class_id(
      class_meta_rsp_fifo_io_in_bits_class_meta_field_type_31_sub_class_id),
    .io_in_bits_class_meta_field_type_32_is_repeated(class_meta_rsp_fifo_io_in_bits_class_meta_field_type_32_is_repeated
      ),
    .io_in_bits_class_meta_field_type_32_field_type(class_meta_rsp_fifo_io_in_bits_class_meta_field_type_32_field_type),
    .io_in_bits_class_meta_field_type_32_sub_class_id(
      class_meta_rsp_fifo_io_in_bits_class_meta_field_type_32_sub_class_id),
    .io_out_ready(class_meta_rsp_fifo_io_out_ready),
    .io_out_valid(class_meta_rsp_fifo_io_out_valid),
    .io_out_bits_class_meta_max_field_num(class_meta_rsp_fifo_io_out_bits_class_meta_max_field_num),
    .io_out_bits_class_meta_field_type_0_is_repeated(class_meta_rsp_fifo_io_out_bits_class_meta_field_type_0_is_repeated
      ),
    .io_out_bits_class_meta_field_type_0_field_type(class_meta_rsp_fifo_io_out_bits_class_meta_field_type_0_field_type),
    .io_out_bits_class_meta_field_type_0_sub_class_id(
      class_meta_rsp_fifo_io_out_bits_class_meta_field_type_0_sub_class_id),
    .io_out_bits_class_meta_field_type_1_is_repeated(class_meta_rsp_fifo_io_out_bits_class_meta_field_type_1_is_repeated
      ),
    .io_out_bits_class_meta_field_type_1_field_type(class_meta_rsp_fifo_io_out_bits_class_meta_field_type_1_field_type),
    .io_out_bits_class_meta_field_type_1_sub_class_id(
      class_meta_rsp_fifo_io_out_bits_class_meta_field_type_1_sub_class_id),
    .io_out_bits_class_meta_field_type_2_is_repeated(class_meta_rsp_fifo_io_out_bits_class_meta_field_type_2_is_repeated
      ),
    .io_out_bits_class_meta_field_type_2_field_type(class_meta_rsp_fifo_io_out_bits_class_meta_field_type_2_field_type),
    .io_out_bits_class_meta_field_type_2_sub_class_id(
      class_meta_rsp_fifo_io_out_bits_class_meta_field_type_2_sub_class_id),
    .io_out_bits_class_meta_field_type_3_is_repeated(class_meta_rsp_fifo_io_out_bits_class_meta_field_type_3_is_repeated
      ),
    .io_out_bits_class_meta_field_type_3_field_type(class_meta_rsp_fifo_io_out_bits_class_meta_field_type_3_field_type),
    .io_out_bits_class_meta_field_type_3_sub_class_id(
      class_meta_rsp_fifo_io_out_bits_class_meta_field_type_3_sub_class_id),
    .io_out_bits_class_meta_field_type_4_is_repeated(class_meta_rsp_fifo_io_out_bits_class_meta_field_type_4_is_repeated
      ),
    .io_out_bits_class_meta_field_type_4_field_type(class_meta_rsp_fifo_io_out_bits_class_meta_field_type_4_field_type),
    .io_out_bits_class_meta_field_type_4_sub_class_id(
      class_meta_rsp_fifo_io_out_bits_class_meta_field_type_4_sub_class_id),
    .io_out_bits_class_meta_field_type_5_is_repeated(class_meta_rsp_fifo_io_out_bits_class_meta_field_type_5_is_repeated
      ),
    .io_out_bits_class_meta_field_type_5_field_type(class_meta_rsp_fifo_io_out_bits_class_meta_field_type_5_field_type),
    .io_out_bits_class_meta_field_type_5_sub_class_id(
      class_meta_rsp_fifo_io_out_bits_class_meta_field_type_5_sub_class_id),
    .io_out_bits_class_meta_field_type_6_is_repeated(class_meta_rsp_fifo_io_out_bits_class_meta_field_type_6_is_repeated
      ),
    .io_out_bits_class_meta_field_type_6_field_type(class_meta_rsp_fifo_io_out_bits_class_meta_field_type_6_field_type),
    .io_out_bits_class_meta_field_type_6_sub_class_id(
      class_meta_rsp_fifo_io_out_bits_class_meta_field_type_6_sub_class_id),
    .io_out_bits_class_meta_field_type_7_is_repeated(class_meta_rsp_fifo_io_out_bits_class_meta_field_type_7_is_repeated
      ),
    .io_out_bits_class_meta_field_type_7_field_type(class_meta_rsp_fifo_io_out_bits_class_meta_field_type_7_field_type),
    .io_out_bits_class_meta_field_type_7_sub_class_id(
      class_meta_rsp_fifo_io_out_bits_class_meta_field_type_7_sub_class_id),
    .io_out_bits_class_meta_field_type_8_is_repeated(class_meta_rsp_fifo_io_out_bits_class_meta_field_type_8_is_repeated
      ),
    .io_out_bits_class_meta_field_type_8_field_type(class_meta_rsp_fifo_io_out_bits_class_meta_field_type_8_field_type),
    .io_out_bits_class_meta_field_type_8_sub_class_id(
      class_meta_rsp_fifo_io_out_bits_class_meta_field_type_8_sub_class_id),
    .io_out_bits_class_meta_field_type_9_is_repeated(class_meta_rsp_fifo_io_out_bits_class_meta_field_type_9_is_repeated
      ),
    .io_out_bits_class_meta_field_type_9_field_type(class_meta_rsp_fifo_io_out_bits_class_meta_field_type_9_field_type),
    .io_out_bits_class_meta_field_type_9_sub_class_id(
      class_meta_rsp_fifo_io_out_bits_class_meta_field_type_9_sub_class_id),
    .io_out_bits_class_meta_field_type_10_is_repeated(
      class_meta_rsp_fifo_io_out_bits_class_meta_field_type_10_is_repeated),
    .io_out_bits_class_meta_field_type_10_field_type(class_meta_rsp_fifo_io_out_bits_class_meta_field_type_10_field_type
      ),
    .io_out_bits_class_meta_field_type_10_sub_class_id(
      class_meta_rsp_fifo_io_out_bits_class_meta_field_type_10_sub_class_id),
    .io_out_bits_class_meta_field_type_11_is_repeated(
      class_meta_rsp_fifo_io_out_bits_class_meta_field_type_11_is_repeated),
    .io_out_bits_class_meta_field_type_11_field_type(class_meta_rsp_fifo_io_out_bits_class_meta_field_type_11_field_type
      ),
    .io_out_bits_class_meta_field_type_11_sub_class_id(
      class_meta_rsp_fifo_io_out_bits_class_meta_field_type_11_sub_class_id),
    .io_out_bits_class_meta_field_type_12_is_repeated(
      class_meta_rsp_fifo_io_out_bits_class_meta_field_type_12_is_repeated),
    .io_out_bits_class_meta_field_type_12_field_type(class_meta_rsp_fifo_io_out_bits_class_meta_field_type_12_field_type
      ),
    .io_out_bits_class_meta_field_type_12_sub_class_id(
      class_meta_rsp_fifo_io_out_bits_class_meta_field_type_12_sub_class_id),
    .io_out_bits_class_meta_field_type_13_is_repeated(
      class_meta_rsp_fifo_io_out_bits_class_meta_field_type_13_is_repeated),
    .io_out_bits_class_meta_field_type_13_field_type(class_meta_rsp_fifo_io_out_bits_class_meta_field_type_13_field_type
      ),
    .io_out_bits_class_meta_field_type_13_sub_class_id(
      class_meta_rsp_fifo_io_out_bits_class_meta_field_type_13_sub_class_id),
    .io_out_bits_class_meta_field_type_14_is_repeated(
      class_meta_rsp_fifo_io_out_bits_class_meta_field_type_14_is_repeated),
    .io_out_bits_class_meta_field_type_14_field_type(class_meta_rsp_fifo_io_out_bits_class_meta_field_type_14_field_type
      ),
    .io_out_bits_class_meta_field_type_14_sub_class_id(
      class_meta_rsp_fifo_io_out_bits_class_meta_field_type_14_sub_class_id),
    .io_out_bits_class_meta_field_type_15_is_repeated(
      class_meta_rsp_fifo_io_out_bits_class_meta_field_type_15_is_repeated),
    .io_out_bits_class_meta_field_type_15_field_type(class_meta_rsp_fifo_io_out_bits_class_meta_field_type_15_field_type
      ),
    .io_out_bits_class_meta_field_type_15_sub_class_id(
      class_meta_rsp_fifo_io_out_bits_class_meta_field_type_15_sub_class_id),
    .io_out_bits_class_meta_field_type_16_is_repeated(
      class_meta_rsp_fifo_io_out_bits_class_meta_field_type_16_is_repeated),
    .io_out_bits_class_meta_field_type_16_field_type(class_meta_rsp_fifo_io_out_bits_class_meta_field_type_16_field_type
      ),
    .io_out_bits_class_meta_field_type_16_sub_class_id(
      class_meta_rsp_fifo_io_out_bits_class_meta_field_type_16_sub_class_id),
    .io_out_bits_class_meta_field_type_17_is_repeated(
      class_meta_rsp_fifo_io_out_bits_class_meta_field_type_17_is_repeated),
    .io_out_bits_class_meta_field_type_17_field_type(class_meta_rsp_fifo_io_out_bits_class_meta_field_type_17_field_type
      ),
    .io_out_bits_class_meta_field_type_17_sub_class_id(
      class_meta_rsp_fifo_io_out_bits_class_meta_field_type_17_sub_class_id),
    .io_out_bits_class_meta_field_type_18_is_repeated(
      class_meta_rsp_fifo_io_out_bits_class_meta_field_type_18_is_repeated),
    .io_out_bits_class_meta_field_type_18_field_type(class_meta_rsp_fifo_io_out_bits_class_meta_field_type_18_field_type
      ),
    .io_out_bits_class_meta_field_type_18_sub_class_id(
      class_meta_rsp_fifo_io_out_bits_class_meta_field_type_18_sub_class_id),
    .io_out_bits_class_meta_field_type_19_is_repeated(
      class_meta_rsp_fifo_io_out_bits_class_meta_field_type_19_is_repeated),
    .io_out_bits_class_meta_field_type_19_field_type(class_meta_rsp_fifo_io_out_bits_class_meta_field_type_19_field_type
      ),
    .io_out_bits_class_meta_field_type_19_sub_class_id(
      class_meta_rsp_fifo_io_out_bits_class_meta_field_type_19_sub_class_id),
    .io_out_bits_class_meta_field_type_20_is_repeated(
      class_meta_rsp_fifo_io_out_bits_class_meta_field_type_20_is_repeated),
    .io_out_bits_class_meta_field_type_20_field_type(class_meta_rsp_fifo_io_out_bits_class_meta_field_type_20_field_type
      ),
    .io_out_bits_class_meta_field_type_20_sub_class_id(
      class_meta_rsp_fifo_io_out_bits_class_meta_field_type_20_sub_class_id),
    .io_out_bits_class_meta_field_type_21_is_repeated(
      class_meta_rsp_fifo_io_out_bits_class_meta_field_type_21_is_repeated),
    .io_out_bits_class_meta_field_type_21_field_type(class_meta_rsp_fifo_io_out_bits_class_meta_field_type_21_field_type
      ),
    .io_out_bits_class_meta_field_type_21_sub_class_id(
      class_meta_rsp_fifo_io_out_bits_class_meta_field_type_21_sub_class_id),
    .io_out_bits_class_meta_field_type_22_is_repeated(
      class_meta_rsp_fifo_io_out_bits_class_meta_field_type_22_is_repeated),
    .io_out_bits_class_meta_field_type_22_field_type(class_meta_rsp_fifo_io_out_bits_class_meta_field_type_22_field_type
      ),
    .io_out_bits_class_meta_field_type_22_sub_class_id(
      class_meta_rsp_fifo_io_out_bits_class_meta_field_type_22_sub_class_id),
    .io_out_bits_class_meta_field_type_23_is_repeated(
      class_meta_rsp_fifo_io_out_bits_class_meta_field_type_23_is_repeated),
    .io_out_bits_class_meta_field_type_23_field_type(class_meta_rsp_fifo_io_out_bits_class_meta_field_type_23_field_type
      ),
    .io_out_bits_class_meta_field_type_23_sub_class_id(
      class_meta_rsp_fifo_io_out_bits_class_meta_field_type_23_sub_class_id),
    .io_out_bits_class_meta_field_type_24_is_repeated(
      class_meta_rsp_fifo_io_out_bits_class_meta_field_type_24_is_repeated),
    .io_out_bits_class_meta_field_type_24_field_type(class_meta_rsp_fifo_io_out_bits_class_meta_field_type_24_field_type
      ),
    .io_out_bits_class_meta_field_type_24_sub_class_id(
      class_meta_rsp_fifo_io_out_bits_class_meta_field_type_24_sub_class_id),
    .io_out_bits_class_meta_field_type_25_is_repeated(
      class_meta_rsp_fifo_io_out_bits_class_meta_field_type_25_is_repeated),
    .io_out_bits_class_meta_field_type_25_field_type(class_meta_rsp_fifo_io_out_bits_class_meta_field_type_25_field_type
      ),
    .io_out_bits_class_meta_field_type_25_sub_class_id(
      class_meta_rsp_fifo_io_out_bits_class_meta_field_type_25_sub_class_id),
    .io_out_bits_class_meta_field_type_26_is_repeated(
      class_meta_rsp_fifo_io_out_bits_class_meta_field_type_26_is_repeated),
    .io_out_bits_class_meta_field_type_26_field_type(class_meta_rsp_fifo_io_out_bits_class_meta_field_type_26_field_type
      ),
    .io_out_bits_class_meta_field_type_26_sub_class_id(
      class_meta_rsp_fifo_io_out_bits_class_meta_field_type_26_sub_class_id),
    .io_out_bits_class_meta_field_type_27_is_repeated(
      class_meta_rsp_fifo_io_out_bits_class_meta_field_type_27_is_repeated),
    .io_out_bits_class_meta_field_type_27_field_type(class_meta_rsp_fifo_io_out_bits_class_meta_field_type_27_field_type
      ),
    .io_out_bits_class_meta_field_type_27_sub_class_id(
      class_meta_rsp_fifo_io_out_bits_class_meta_field_type_27_sub_class_id),
    .io_out_bits_class_meta_field_type_28_is_repeated(
      class_meta_rsp_fifo_io_out_bits_class_meta_field_type_28_is_repeated),
    .io_out_bits_class_meta_field_type_28_field_type(class_meta_rsp_fifo_io_out_bits_class_meta_field_type_28_field_type
      ),
    .io_out_bits_class_meta_field_type_28_sub_class_id(
      class_meta_rsp_fifo_io_out_bits_class_meta_field_type_28_sub_class_id),
    .io_out_bits_class_meta_field_type_29_is_repeated(
      class_meta_rsp_fifo_io_out_bits_class_meta_field_type_29_is_repeated),
    .io_out_bits_class_meta_field_type_29_field_type(class_meta_rsp_fifo_io_out_bits_class_meta_field_type_29_field_type
      ),
    .io_out_bits_class_meta_field_type_29_sub_class_id(
      class_meta_rsp_fifo_io_out_bits_class_meta_field_type_29_sub_class_id),
    .io_out_bits_class_meta_field_type_30_is_repeated(
      class_meta_rsp_fifo_io_out_bits_class_meta_field_type_30_is_repeated),
    .io_out_bits_class_meta_field_type_30_field_type(class_meta_rsp_fifo_io_out_bits_class_meta_field_type_30_field_type
      ),
    .io_out_bits_class_meta_field_type_30_sub_class_id(
      class_meta_rsp_fifo_io_out_bits_class_meta_field_type_30_sub_class_id),
    .io_out_bits_class_meta_field_type_31_is_repeated(
      class_meta_rsp_fifo_io_out_bits_class_meta_field_type_31_is_repeated),
    .io_out_bits_class_meta_field_type_31_field_type(class_meta_rsp_fifo_io_out_bits_class_meta_field_type_31_field_type
      ),
    .io_out_bits_class_meta_field_type_31_sub_class_id(
      class_meta_rsp_fifo_io_out_bits_class_meta_field_type_31_sub_class_id),
    .io_out_bits_class_meta_field_type_32_is_repeated(
      class_meta_rsp_fifo_io_out_bits_class_meta_field_type_32_is_repeated),
    .io_out_bits_class_meta_field_type_32_field_type(class_meta_rsp_fifo_io_out_bits_class_meta_field_type_32_field_type
      ),
    .io_out_bits_class_meta_field_type_32_sub_class_id(
      class_meta_rsp_fifo_io_out_bits_class_meta_field_type_32_sub_class_id)
  );
  assign io_meta_in_ready = meta_in_fifo_io_in_ready; // @[Serializerhw.scala 35:41]
  assign io_host_data_in_ready = 1'h1; // @[Serializerhw.scala 36:41]
  assign io_host_data_cmd_valid = _T_4 ? 1'h0 : _GEN_8578; // @[Conditional.scala 40:58 Util.scala 13:25]
  assign io_host_data_cmd_bits_vaddr = _T_4 ? 64'h0 : _GEN_8579; // @[Conditional.scala 40:58 Util.scala 13:25]
  assign io_host_data_cmd_bits_length = _T_4 ? 32'h0 : _GEN_8580; // @[Conditional.scala 40:58 Util.scala 13:25]
  assign io_class_meta_req_valid = _T_4 ? _T_5 : _GEN_8587; // @[Conditional.scala 40:58]
  assign io_class_meta_req_bits_class_id = _GEN_8601[9:0];
  assign io_done_valid = _T_4 ? 1'h0 : _GEN_8591; // @[Conditional.scala 40:58 Util.scala 13:25]
  assign counter_3_0 = counter_3;
  assign counter_2_0 = counter_2;
  assign counter_8 = counter;
  assign counter_1_1 = counter_1;
  assign meta_in_fifo_clock = clock;
  assign meta_in_fifo_reset = reset;
  assign meta_in_fifo_io_in_valid = io_meta_in_valid; // @[Serializerhw.scala 35:41]
  assign meta_in_fifo_io_in_bits_class_id = io_meta_in_bits_class_id; // @[Serializerhw.scala 35:41]
  assign meta_in_fifo_io_in_bits_host_base_addr = io_meta_in_bits_host_base_addr; // @[Serializerhw.scala 35:41]
  assign meta_in_fifo_io_out_ready = state == 5'h6 & io_class_meta_req_ready; // @[Serializerhw.scala 89:68]
  assign class_meta_rsp_fifo_clock = clock;
  assign class_meta_rsp_fifo_reset = reset;
  assign class_meta_rsp_fifo_io_in_valid = io_class_meta_rsp_valid; // @[Serializerhw.scala 37:41]
  assign class_meta_rsp_fifo_io_in_bits_class_meta_max_field_num = io_class_meta_rsp_bits_class_meta_max_field_num; // @[Serializerhw.scala 37:41]
  assign class_meta_rsp_fifo_io_in_bits_class_meta_field_type_0_is_repeated =
    io_class_meta_rsp_bits_class_meta_field_type_0_is_repeated; // @[Serializerhw.scala 37:41]
  assign class_meta_rsp_fifo_io_in_bits_class_meta_field_type_0_field_type =
    io_class_meta_rsp_bits_class_meta_field_type_0_field_type; // @[Serializerhw.scala 37:41]
  assign class_meta_rsp_fifo_io_in_bits_class_meta_field_type_0_sub_class_id =
    io_class_meta_rsp_bits_class_meta_field_type_0_sub_class_id; // @[Serializerhw.scala 37:41]
  assign class_meta_rsp_fifo_io_in_bits_class_meta_field_type_1_is_repeated =
    io_class_meta_rsp_bits_class_meta_field_type_1_is_repeated; // @[Serializerhw.scala 37:41]
  assign class_meta_rsp_fifo_io_in_bits_class_meta_field_type_1_field_type =
    io_class_meta_rsp_bits_class_meta_field_type_1_field_type; // @[Serializerhw.scala 37:41]
  assign class_meta_rsp_fifo_io_in_bits_class_meta_field_type_1_sub_class_id =
    io_class_meta_rsp_bits_class_meta_field_type_1_sub_class_id; // @[Serializerhw.scala 37:41]
  assign class_meta_rsp_fifo_io_in_bits_class_meta_field_type_2_is_repeated =
    io_class_meta_rsp_bits_class_meta_field_type_2_is_repeated; // @[Serializerhw.scala 37:41]
  assign class_meta_rsp_fifo_io_in_bits_class_meta_field_type_2_field_type =
    io_class_meta_rsp_bits_class_meta_field_type_2_field_type; // @[Serializerhw.scala 37:41]
  assign class_meta_rsp_fifo_io_in_bits_class_meta_field_type_2_sub_class_id =
    io_class_meta_rsp_bits_class_meta_field_type_2_sub_class_id; // @[Serializerhw.scala 37:41]
  assign class_meta_rsp_fifo_io_in_bits_class_meta_field_type_3_is_repeated =
    io_class_meta_rsp_bits_class_meta_field_type_3_is_repeated; // @[Serializerhw.scala 37:41]
  assign class_meta_rsp_fifo_io_in_bits_class_meta_field_type_3_field_type =
    io_class_meta_rsp_bits_class_meta_field_type_3_field_type; // @[Serializerhw.scala 37:41]
  assign class_meta_rsp_fifo_io_in_bits_class_meta_field_type_3_sub_class_id =
    io_class_meta_rsp_bits_class_meta_field_type_3_sub_class_id; // @[Serializerhw.scala 37:41]
  assign class_meta_rsp_fifo_io_in_bits_class_meta_field_type_4_is_repeated =
    io_class_meta_rsp_bits_class_meta_field_type_4_is_repeated; // @[Serializerhw.scala 37:41]
  assign class_meta_rsp_fifo_io_in_bits_class_meta_field_type_4_field_type =
    io_class_meta_rsp_bits_class_meta_field_type_4_field_type; // @[Serializerhw.scala 37:41]
  assign class_meta_rsp_fifo_io_in_bits_class_meta_field_type_4_sub_class_id =
    io_class_meta_rsp_bits_class_meta_field_type_4_sub_class_id; // @[Serializerhw.scala 37:41]
  assign class_meta_rsp_fifo_io_in_bits_class_meta_field_type_5_is_repeated =
    io_class_meta_rsp_bits_class_meta_field_type_5_is_repeated; // @[Serializerhw.scala 37:41]
  assign class_meta_rsp_fifo_io_in_bits_class_meta_field_type_5_field_type =
    io_class_meta_rsp_bits_class_meta_field_type_5_field_type; // @[Serializerhw.scala 37:41]
  assign class_meta_rsp_fifo_io_in_bits_class_meta_field_type_5_sub_class_id =
    io_class_meta_rsp_bits_class_meta_field_type_5_sub_class_id; // @[Serializerhw.scala 37:41]
  assign class_meta_rsp_fifo_io_in_bits_class_meta_field_type_6_is_repeated =
    io_class_meta_rsp_bits_class_meta_field_type_6_is_repeated; // @[Serializerhw.scala 37:41]
  assign class_meta_rsp_fifo_io_in_bits_class_meta_field_type_6_field_type =
    io_class_meta_rsp_bits_class_meta_field_type_6_field_type; // @[Serializerhw.scala 37:41]
  assign class_meta_rsp_fifo_io_in_bits_class_meta_field_type_6_sub_class_id =
    io_class_meta_rsp_bits_class_meta_field_type_6_sub_class_id; // @[Serializerhw.scala 37:41]
  assign class_meta_rsp_fifo_io_in_bits_class_meta_field_type_7_is_repeated =
    io_class_meta_rsp_bits_class_meta_field_type_7_is_repeated; // @[Serializerhw.scala 37:41]
  assign class_meta_rsp_fifo_io_in_bits_class_meta_field_type_7_field_type =
    io_class_meta_rsp_bits_class_meta_field_type_7_field_type; // @[Serializerhw.scala 37:41]
  assign class_meta_rsp_fifo_io_in_bits_class_meta_field_type_7_sub_class_id =
    io_class_meta_rsp_bits_class_meta_field_type_7_sub_class_id; // @[Serializerhw.scala 37:41]
  assign class_meta_rsp_fifo_io_in_bits_class_meta_field_type_8_is_repeated =
    io_class_meta_rsp_bits_class_meta_field_type_8_is_repeated; // @[Serializerhw.scala 37:41]
  assign class_meta_rsp_fifo_io_in_bits_class_meta_field_type_8_field_type =
    io_class_meta_rsp_bits_class_meta_field_type_8_field_type; // @[Serializerhw.scala 37:41]
  assign class_meta_rsp_fifo_io_in_bits_class_meta_field_type_8_sub_class_id =
    io_class_meta_rsp_bits_class_meta_field_type_8_sub_class_id; // @[Serializerhw.scala 37:41]
  assign class_meta_rsp_fifo_io_in_bits_class_meta_field_type_9_is_repeated =
    io_class_meta_rsp_bits_class_meta_field_type_9_is_repeated; // @[Serializerhw.scala 37:41]
  assign class_meta_rsp_fifo_io_in_bits_class_meta_field_type_9_field_type =
    io_class_meta_rsp_bits_class_meta_field_type_9_field_type; // @[Serializerhw.scala 37:41]
  assign class_meta_rsp_fifo_io_in_bits_class_meta_field_type_9_sub_class_id =
    io_class_meta_rsp_bits_class_meta_field_type_9_sub_class_id; // @[Serializerhw.scala 37:41]
  assign class_meta_rsp_fifo_io_in_bits_class_meta_field_type_10_is_repeated =
    io_class_meta_rsp_bits_class_meta_field_type_10_is_repeated; // @[Serializerhw.scala 37:41]
  assign class_meta_rsp_fifo_io_in_bits_class_meta_field_type_10_field_type =
    io_class_meta_rsp_bits_class_meta_field_type_10_field_type; // @[Serializerhw.scala 37:41]
  assign class_meta_rsp_fifo_io_in_bits_class_meta_field_type_10_sub_class_id =
    io_class_meta_rsp_bits_class_meta_field_type_10_sub_class_id; // @[Serializerhw.scala 37:41]
  assign class_meta_rsp_fifo_io_in_bits_class_meta_field_type_11_is_repeated =
    io_class_meta_rsp_bits_class_meta_field_type_11_is_repeated; // @[Serializerhw.scala 37:41]
  assign class_meta_rsp_fifo_io_in_bits_class_meta_field_type_11_field_type =
    io_class_meta_rsp_bits_class_meta_field_type_11_field_type; // @[Serializerhw.scala 37:41]
  assign class_meta_rsp_fifo_io_in_bits_class_meta_field_type_11_sub_class_id =
    io_class_meta_rsp_bits_class_meta_field_type_11_sub_class_id; // @[Serializerhw.scala 37:41]
  assign class_meta_rsp_fifo_io_in_bits_class_meta_field_type_12_is_repeated =
    io_class_meta_rsp_bits_class_meta_field_type_12_is_repeated; // @[Serializerhw.scala 37:41]
  assign class_meta_rsp_fifo_io_in_bits_class_meta_field_type_12_field_type =
    io_class_meta_rsp_bits_class_meta_field_type_12_field_type; // @[Serializerhw.scala 37:41]
  assign class_meta_rsp_fifo_io_in_bits_class_meta_field_type_12_sub_class_id =
    io_class_meta_rsp_bits_class_meta_field_type_12_sub_class_id; // @[Serializerhw.scala 37:41]
  assign class_meta_rsp_fifo_io_in_bits_class_meta_field_type_13_is_repeated =
    io_class_meta_rsp_bits_class_meta_field_type_13_is_repeated; // @[Serializerhw.scala 37:41]
  assign class_meta_rsp_fifo_io_in_bits_class_meta_field_type_13_field_type =
    io_class_meta_rsp_bits_class_meta_field_type_13_field_type; // @[Serializerhw.scala 37:41]
  assign class_meta_rsp_fifo_io_in_bits_class_meta_field_type_13_sub_class_id =
    io_class_meta_rsp_bits_class_meta_field_type_13_sub_class_id; // @[Serializerhw.scala 37:41]
  assign class_meta_rsp_fifo_io_in_bits_class_meta_field_type_14_is_repeated =
    io_class_meta_rsp_bits_class_meta_field_type_14_is_repeated; // @[Serializerhw.scala 37:41]
  assign class_meta_rsp_fifo_io_in_bits_class_meta_field_type_14_field_type =
    io_class_meta_rsp_bits_class_meta_field_type_14_field_type; // @[Serializerhw.scala 37:41]
  assign class_meta_rsp_fifo_io_in_bits_class_meta_field_type_14_sub_class_id =
    io_class_meta_rsp_bits_class_meta_field_type_14_sub_class_id; // @[Serializerhw.scala 37:41]
  assign class_meta_rsp_fifo_io_in_bits_class_meta_field_type_15_is_repeated =
    io_class_meta_rsp_bits_class_meta_field_type_15_is_repeated; // @[Serializerhw.scala 37:41]
  assign class_meta_rsp_fifo_io_in_bits_class_meta_field_type_15_field_type =
    io_class_meta_rsp_bits_class_meta_field_type_15_field_type; // @[Serializerhw.scala 37:41]
  assign class_meta_rsp_fifo_io_in_bits_class_meta_field_type_15_sub_class_id =
    io_class_meta_rsp_bits_class_meta_field_type_15_sub_class_id; // @[Serializerhw.scala 37:41]
  assign class_meta_rsp_fifo_io_in_bits_class_meta_field_type_16_is_repeated =
    io_class_meta_rsp_bits_class_meta_field_type_16_is_repeated; // @[Serializerhw.scala 37:41]
  assign class_meta_rsp_fifo_io_in_bits_class_meta_field_type_16_field_type =
    io_class_meta_rsp_bits_class_meta_field_type_16_field_type; // @[Serializerhw.scala 37:41]
  assign class_meta_rsp_fifo_io_in_bits_class_meta_field_type_16_sub_class_id =
    io_class_meta_rsp_bits_class_meta_field_type_16_sub_class_id; // @[Serializerhw.scala 37:41]
  assign class_meta_rsp_fifo_io_in_bits_class_meta_field_type_17_is_repeated =
    io_class_meta_rsp_bits_class_meta_field_type_17_is_repeated; // @[Serializerhw.scala 37:41]
  assign class_meta_rsp_fifo_io_in_bits_class_meta_field_type_17_field_type =
    io_class_meta_rsp_bits_class_meta_field_type_17_field_type; // @[Serializerhw.scala 37:41]
  assign class_meta_rsp_fifo_io_in_bits_class_meta_field_type_17_sub_class_id =
    io_class_meta_rsp_bits_class_meta_field_type_17_sub_class_id; // @[Serializerhw.scala 37:41]
  assign class_meta_rsp_fifo_io_in_bits_class_meta_field_type_18_is_repeated =
    io_class_meta_rsp_bits_class_meta_field_type_18_is_repeated; // @[Serializerhw.scala 37:41]
  assign class_meta_rsp_fifo_io_in_bits_class_meta_field_type_18_field_type =
    io_class_meta_rsp_bits_class_meta_field_type_18_field_type; // @[Serializerhw.scala 37:41]
  assign class_meta_rsp_fifo_io_in_bits_class_meta_field_type_18_sub_class_id =
    io_class_meta_rsp_bits_class_meta_field_type_18_sub_class_id; // @[Serializerhw.scala 37:41]
  assign class_meta_rsp_fifo_io_in_bits_class_meta_field_type_19_is_repeated =
    io_class_meta_rsp_bits_class_meta_field_type_19_is_repeated; // @[Serializerhw.scala 37:41]
  assign class_meta_rsp_fifo_io_in_bits_class_meta_field_type_19_field_type =
    io_class_meta_rsp_bits_class_meta_field_type_19_field_type; // @[Serializerhw.scala 37:41]
  assign class_meta_rsp_fifo_io_in_bits_class_meta_field_type_19_sub_class_id =
    io_class_meta_rsp_bits_class_meta_field_type_19_sub_class_id; // @[Serializerhw.scala 37:41]
  assign class_meta_rsp_fifo_io_in_bits_class_meta_field_type_20_is_repeated =
    io_class_meta_rsp_bits_class_meta_field_type_20_is_repeated; // @[Serializerhw.scala 37:41]
  assign class_meta_rsp_fifo_io_in_bits_class_meta_field_type_20_field_type =
    io_class_meta_rsp_bits_class_meta_field_type_20_field_type; // @[Serializerhw.scala 37:41]
  assign class_meta_rsp_fifo_io_in_bits_class_meta_field_type_20_sub_class_id =
    io_class_meta_rsp_bits_class_meta_field_type_20_sub_class_id; // @[Serializerhw.scala 37:41]
  assign class_meta_rsp_fifo_io_in_bits_class_meta_field_type_21_is_repeated =
    io_class_meta_rsp_bits_class_meta_field_type_21_is_repeated; // @[Serializerhw.scala 37:41]
  assign class_meta_rsp_fifo_io_in_bits_class_meta_field_type_21_field_type =
    io_class_meta_rsp_bits_class_meta_field_type_21_field_type; // @[Serializerhw.scala 37:41]
  assign class_meta_rsp_fifo_io_in_bits_class_meta_field_type_21_sub_class_id =
    io_class_meta_rsp_bits_class_meta_field_type_21_sub_class_id; // @[Serializerhw.scala 37:41]
  assign class_meta_rsp_fifo_io_in_bits_class_meta_field_type_22_is_repeated =
    io_class_meta_rsp_bits_class_meta_field_type_22_is_repeated; // @[Serializerhw.scala 37:41]
  assign class_meta_rsp_fifo_io_in_bits_class_meta_field_type_22_field_type =
    io_class_meta_rsp_bits_class_meta_field_type_22_field_type; // @[Serializerhw.scala 37:41]
  assign class_meta_rsp_fifo_io_in_bits_class_meta_field_type_22_sub_class_id =
    io_class_meta_rsp_bits_class_meta_field_type_22_sub_class_id; // @[Serializerhw.scala 37:41]
  assign class_meta_rsp_fifo_io_in_bits_class_meta_field_type_23_is_repeated =
    io_class_meta_rsp_bits_class_meta_field_type_23_is_repeated; // @[Serializerhw.scala 37:41]
  assign class_meta_rsp_fifo_io_in_bits_class_meta_field_type_23_field_type =
    io_class_meta_rsp_bits_class_meta_field_type_23_field_type; // @[Serializerhw.scala 37:41]
  assign class_meta_rsp_fifo_io_in_bits_class_meta_field_type_23_sub_class_id =
    io_class_meta_rsp_bits_class_meta_field_type_23_sub_class_id; // @[Serializerhw.scala 37:41]
  assign class_meta_rsp_fifo_io_in_bits_class_meta_field_type_24_is_repeated =
    io_class_meta_rsp_bits_class_meta_field_type_24_is_repeated; // @[Serializerhw.scala 37:41]
  assign class_meta_rsp_fifo_io_in_bits_class_meta_field_type_24_field_type =
    io_class_meta_rsp_bits_class_meta_field_type_24_field_type; // @[Serializerhw.scala 37:41]
  assign class_meta_rsp_fifo_io_in_bits_class_meta_field_type_24_sub_class_id =
    io_class_meta_rsp_bits_class_meta_field_type_24_sub_class_id; // @[Serializerhw.scala 37:41]
  assign class_meta_rsp_fifo_io_in_bits_class_meta_field_type_25_is_repeated =
    io_class_meta_rsp_bits_class_meta_field_type_25_is_repeated; // @[Serializerhw.scala 37:41]
  assign class_meta_rsp_fifo_io_in_bits_class_meta_field_type_25_field_type =
    io_class_meta_rsp_bits_class_meta_field_type_25_field_type; // @[Serializerhw.scala 37:41]
  assign class_meta_rsp_fifo_io_in_bits_class_meta_field_type_25_sub_class_id =
    io_class_meta_rsp_bits_class_meta_field_type_25_sub_class_id; // @[Serializerhw.scala 37:41]
  assign class_meta_rsp_fifo_io_in_bits_class_meta_field_type_26_is_repeated =
    io_class_meta_rsp_bits_class_meta_field_type_26_is_repeated; // @[Serializerhw.scala 37:41]
  assign class_meta_rsp_fifo_io_in_bits_class_meta_field_type_26_field_type =
    io_class_meta_rsp_bits_class_meta_field_type_26_field_type; // @[Serializerhw.scala 37:41]
  assign class_meta_rsp_fifo_io_in_bits_class_meta_field_type_26_sub_class_id =
    io_class_meta_rsp_bits_class_meta_field_type_26_sub_class_id; // @[Serializerhw.scala 37:41]
  assign class_meta_rsp_fifo_io_in_bits_class_meta_field_type_27_is_repeated =
    io_class_meta_rsp_bits_class_meta_field_type_27_is_repeated; // @[Serializerhw.scala 37:41]
  assign class_meta_rsp_fifo_io_in_bits_class_meta_field_type_27_field_type =
    io_class_meta_rsp_bits_class_meta_field_type_27_field_type; // @[Serializerhw.scala 37:41]
  assign class_meta_rsp_fifo_io_in_bits_class_meta_field_type_27_sub_class_id =
    io_class_meta_rsp_bits_class_meta_field_type_27_sub_class_id; // @[Serializerhw.scala 37:41]
  assign class_meta_rsp_fifo_io_in_bits_class_meta_field_type_28_is_repeated =
    io_class_meta_rsp_bits_class_meta_field_type_28_is_repeated; // @[Serializerhw.scala 37:41]
  assign class_meta_rsp_fifo_io_in_bits_class_meta_field_type_28_field_type =
    io_class_meta_rsp_bits_class_meta_field_type_28_field_type; // @[Serializerhw.scala 37:41]
  assign class_meta_rsp_fifo_io_in_bits_class_meta_field_type_28_sub_class_id =
    io_class_meta_rsp_bits_class_meta_field_type_28_sub_class_id; // @[Serializerhw.scala 37:41]
  assign class_meta_rsp_fifo_io_in_bits_class_meta_field_type_29_is_repeated =
    io_class_meta_rsp_bits_class_meta_field_type_29_is_repeated; // @[Serializerhw.scala 37:41]
  assign class_meta_rsp_fifo_io_in_bits_class_meta_field_type_29_field_type =
    io_class_meta_rsp_bits_class_meta_field_type_29_field_type; // @[Serializerhw.scala 37:41]
  assign class_meta_rsp_fifo_io_in_bits_class_meta_field_type_29_sub_class_id =
    io_class_meta_rsp_bits_class_meta_field_type_29_sub_class_id; // @[Serializerhw.scala 37:41]
  assign class_meta_rsp_fifo_io_in_bits_class_meta_field_type_30_is_repeated =
    io_class_meta_rsp_bits_class_meta_field_type_30_is_repeated; // @[Serializerhw.scala 37:41]
  assign class_meta_rsp_fifo_io_in_bits_class_meta_field_type_30_field_type =
    io_class_meta_rsp_bits_class_meta_field_type_30_field_type; // @[Serializerhw.scala 37:41]
  assign class_meta_rsp_fifo_io_in_bits_class_meta_field_type_30_sub_class_id =
    io_class_meta_rsp_bits_class_meta_field_type_30_sub_class_id; // @[Serializerhw.scala 37:41]
  assign class_meta_rsp_fifo_io_in_bits_class_meta_field_type_31_is_repeated =
    io_class_meta_rsp_bits_class_meta_field_type_31_is_repeated; // @[Serializerhw.scala 37:41]
  assign class_meta_rsp_fifo_io_in_bits_class_meta_field_type_31_field_type =
    io_class_meta_rsp_bits_class_meta_field_type_31_field_type; // @[Serializerhw.scala 37:41]
  assign class_meta_rsp_fifo_io_in_bits_class_meta_field_type_31_sub_class_id =
    io_class_meta_rsp_bits_class_meta_field_type_31_sub_class_id; // @[Serializerhw.scala 37:41]
  assign class_meta_rsp_fifo_io_in_bits_class_meta_field_type_32_is_repeated =
    io_class_meta_rsp_bits_class_meta_field_type_32_is_repeated; // @[Serializerhw.scala 37:41]
  assign class_meta_rsp_fifo_io_in_bits_class_meta_field_type_32_field_type =
    io_class_meta_rsp_bits_class_meta_field_type_32_field_type; // @[Serializerhw.scala 37:41]
  assign class_meta_rsp_fifo_io_in_bits_class_meta_field_type_32_sub_class_id =
    io_class_meta_rsp_bits_class_meta_field_type_32_sub_class_id; // @[Serializerhw.scala 37:41]
  assign class_meta_rsp_fifo_io_out_ready = state == 5'h11; // @[Serializerhw.scala 90:54]
  always @(posedge clock) begin
    if (reset) begin // @[Collector.scala 169:42]
      counter <= 32'h0; // @[Collector.scala 169:42]
    end else if (_T) begin // @[Collector.scala 170:34]
      counter <= _counter_T_1; // @[Collector.scala 171:41]
    end
    if (reset) begin // @[Collector.scala 169:42]
      counter_1 <= 32'h0; // @[Collector.scala 169:42]
    end else if (_T_1) begin // @[Collector.scala 170:34]
      counter_1 <= _counter_T_3; // @[Collector.scala 171:41]
    end
    if (reset) begin // @[Collector.scala 169:42]
      counter_2 <= 32'h0; // @[Collector.scala 169:42]
    end else if (_T_2) begin // @[Collector.scala 170:34]
      counter_2 <= _counter_T_5; // @[Collector.scala 171:41]
    end
    if (reset) begin // @[Collector.scala 169:42]
      counter_3 <= 32'h0; // @[Collector.scala 169:42]
    end else if (io_done_valid) begin // @[Collector.scala 170:34]
      counter_3 <= _counter_T_7; // @[Collector.scala 171:41]
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h0 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_0_field_type_0_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_0_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h0 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_0_field_type_0_field_type <= _field_stack_stack_num_field_type_0_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h0 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_0_field_type_0_sub_class_id <= _field_stack_stack_num_field_type_0_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h0 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_0_field_type_1_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_1_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h0 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_0_field_type_1_field_type <= _field_stack_stack_num_field_type_1_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h0 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_0_field_type_1_sub_class_id <= _field_stack_stack_num_field_type_1_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h0 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_0_field_type_2_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_2_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h0 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_0_field_type_2_field_type <= _field_stack_stack_num_field_type_2_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h0 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_0_field_type_2_sub_class_id <= _field_stack_stack_num_field_type_2_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h0 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_0_field_type_3_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_3_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h0 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_0_field_type_3_field_type <= _field_stack_stack_num_field_type_3_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h0 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_0_field_type_3_sub_class_id <= _field_stack_stack_num_field_type_3_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h0 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_0_field_type_4_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_4_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h0 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_0_field_type_4_field_type <= _field_stack_stack_num_field_type_4_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h0 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_0_field_type_4_sub_class_id <= _field_stack_stack_num_field_type_4_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h0 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_0_field_type_5_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_5_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h0 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_0_field_type_5_field_type <= _field_stack_stack_num_field_type_5_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h0 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_0_field_type_5_sub_class_id <= _field_stack_stack_num_field_type_5_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h0 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_0_field_type_6_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_6_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h0 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_0_field_type_6_field_type <= _field_stack_stack_num_field_type_6_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h0 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_0_field_type_6_sub_class_id <= _field_stack_stack_num_field_type_6_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h0 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_0_field_type_7_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_7_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h0 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_0_field_type_7_field_type <= _field_stack_stack_num_field_type_7_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h0 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_0_field_type_7_sub_class_id <= _field_stack_stack_num_field_type_7_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h0 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_0_field_type_8_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_8_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h0 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_0_field_type_8_field_type <= _field_stack_stack_num_field_type_8_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h0 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_0_field_type_8_sub_class_id <= _field_stack_stack_num_field_type_8_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h0 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_0_field_type_9_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_9_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h0 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_0_field_type_9_field_type <= _field_stack_stack_num_field_type_9_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h0 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_0_field_type_9_sub_class_id <= _field_stack_stack_num_field_type_9_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h0 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_0_field_type_10_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_10_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h0 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_0_field_type_10_field_type <= _field_stack_stack_num_field_type_10_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h0 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_0_field_type_10_sub_class_id <= _field_stack_stack_num_field_type_10_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h0 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_0_field_type_11_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_11_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h0 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_0_field_type_11_field_type <= _field_stack_stack_num_field_type_11_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h0 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_0_field_type_11_sub_class_id <= _field_stack_stack_num_field_type_11_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h0 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_0_field_type_12_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_12_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h0 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_0_field_type_12_field_type <= _field_stack_stack_num_field_type_12_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h0 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_0_field_type_12_sub_class_id <= _field_stack_stack_num_field_type_12_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h0 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_0_field_type_13_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_13_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h0 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_0_field_type_13_field_type <= _field_stack_stack_num_field_type_13_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h0 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_0_field_type_13_sub_class_id <= _field_stack_stack_num_field_type_13_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h0 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_0_field_type_14_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_14_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h0 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_0_field_type_14_field_type <= _field_stack_stack_num_field_type_14_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h0 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_0_field_type_14_sub_class_id <= _field_stack_stack_num_field_type_14_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h0 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_0_field_type_15_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_15_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h0 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_0_field_type_15_field_type <= _field_stack_stack_num_field_type_15_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h0 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_0_field_type_15_sub_class_id <= _field_stack_stack_num_field_type_15_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h0 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_0_field_type_16_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_16_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h0 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_0_field_type_16_field_type <= _field_stack_stack_num_field_type_16_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h0 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_0_field_type_16_sub_class_id <= _field_stack_stack_num_field_type_16_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h0 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_0_field_type_17_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_17_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h0 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_0_field_type_17_field_type <= _field_stack_stack_num_field_type_17_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h0 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_0_field_type_17_sub_class_id <= _field_stack_stack_num_field_type_17_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h0 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_0_field_type_18_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_18_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h0 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_0_field_type_18_field_type <= _field_stack_stack_num_field_type_18_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h0 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_0_field_type_18_sub_class_id <= _field_stack_stack_num_field_type_18_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h0 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_0_field_type_19_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_19_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h0 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_0_field_type_19_field_type <= _field_stack_stack_num_field_type_19_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h0 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_0_field_type_19_sub_class_id <= _field_stack_stack_num_field_type_19_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h0 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_0_field_type_20_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_20_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h0 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_0_field_type_20_field_type <= _field_stack_stack_num_field_type_20_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h0 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_0_field_type_20_sub_class_id <= _field_stack_stack_num_field_type_20_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h0 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_0_field_type_21_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_21_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h0 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_0_field_type_21_field_type <= _field_stack_stack_num_field_type_21_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h0 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_0_field_type_21_sub_class_id <= _field_stack_stack_num_field_type_21_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h0 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_0_field_type_22_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_22_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h0 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_0_field_type_22_field_type <= _field_stack_stack_num_field_type_22_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h0 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_0_field_type_22_sub_class_id <= _field_stack_stack_num_field_type_22_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h0 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_0_field_type_23_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_23_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h0 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_0_field_type_23_field_type <= _field_stack_stack_num_field_type_23_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h0 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_0_field_type_23_sub_class_id <= _field_stack_stack_num_field_type_23_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h0 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_0_field_type_24_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_24_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h0 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_0_field_type_24_field_type <= _field_stack_stack_num_field_type_24_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h0 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_0_field_type_24_sub_class_id <= _field_stack_stack_num_field_type_24_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h0 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_0_field_type_25_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_25_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h0 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_0_field_type_25_field_type <= _field_stack_stack_num_field_type_25_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h0 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_0_field_type_25_sub_class_id <= _field_stack_stack_num_field_type_25_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h0 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_0_field_type_26_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_26_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h0 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_0_field_type_26_field_type <= _field_stack_stack_num_field_type_26_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h0 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_0_field_type_26_sub_class_id <= _field_stack_stack_num_field_type_26_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h0 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_0_field_type_27_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_27_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h0 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_0_field_type_27_field_type <= _field_stack_stack_num_field_type_27_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h0 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_0_field_type_27_sub_class_id <= _field_stack_stack_num_field_type_27_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h0 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_0_field_type_28_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_28_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h0 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_0_field_type_28_field_type <= _field_stack_stack_num_field_type_28_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h0 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_0_field_type_28_sub_class_id <= _field_stack_stack_num_field_type_28_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h0 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_0_field_type_29_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_29_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h0 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_0_field_type_29_field_type <= _field_stack_stack_num_field_type_29_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h0 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_0_field_type_29_sub_class_id <= _field_stack_stack_num_field_type_29_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h0 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_0_field_type_30_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_30_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h0 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_0_field_type_30_field_type <= _field_stack_stack_num_field_type_30_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h0 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_0_field_type_30_sub_class_id <= _field_stack_stack_num_field_type_30_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h0 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_0_field_type_31_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_31_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h0 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_0_field_type_31_field_type <= _field_stack_stack_num_field_type_31_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h0 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_0_field_type_31_sub_class_id <= _field_stack_stack_num_field_type_31_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h0 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_0_field_type_32_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_32_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h0 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_0_field_type_32_field_type <= _field_stack_stack_num_field_type_32_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h0 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_0_field_type_32_sub_class_id <= _field_stack_stack_num_field_type_32_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h1 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_1_field_type_0_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_0_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h1 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_1_field_type_0_field_type <= _field_stack_stack_num_field_type_0_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h1 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_1_field_type_0_sub_class_id <= _field_stack_stack_num_field_type_0_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h1 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_1_field_type_1_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_1_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h1 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_1_field_type_1_field_type <= _field_stack_stack_num_field_type_1_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h1 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_1_field_type_1_sub_class_id <= _field_stack_stack_num_field_type_1_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h1 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_1_field_type_2_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_2_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h1 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_1_field_type_2_field_type <= _field_stack_stack_num_field_type_2_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h1 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_1_field_type_2_sub_class_id <= _field_stack_stack_num_field_type_2_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h1 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_1_field_type_3_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_3_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h1 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_1_field_type_3_field_type <= _field_stack_stack_num_field_type_3_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h1 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_1_field_type_3_sub_class_id <= _field_stack_stack_num_field_type_3_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h1 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_1_field_type_4_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_4_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h1 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_1_field_type_4_field_type <= _field_stack_stack_num_field_type_4_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h1 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_1_field_type_4_sub_class_id <= _field_stack_stack_num_field_type_4_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h1 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_1_field_type_5_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_5_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h1 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_1_field_type_5_field_type <= _field_stack_stack_num_field_type_5_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h1 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_1_field_type_5_sub_class_id <= _field_stack_stack_num_field_type_5_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h1 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_1_field_type_6_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_6_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h1 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_1_field_type_6_field_type <= _field_stack_stack_num_field_type_6_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h1 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_1_field_type_6_sub_class_id <= _field_stack_stack_num_field_type_6_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h1 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_1_field_type_7_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_7_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h1 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_1_field_type_7_field_type <= _field_stack_stack_num_field_type_7_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h1 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_1_field_type_7_sub_class_id <= _field_stack_stack_num_field_type_7_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h1 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_1_field_type_8_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_8_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h1 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_1_field_type_8_field_type <= _field_stack_stack_num_field_type_8_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h1 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_1_field_type_8_sub_class_id <= _field_stack_stack_num_field_type_8_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h1 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_1_field_type_9_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_9_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h1 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_1_field_type_9_field_type <= _field_stack_stack_num_field_type_9_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h1 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_1_field_type_9_sub_class_id <= _field_stack_stack_num_field_type_9_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h1 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_1_field_type_10_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_10_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h1 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_1_field_type_10_field_type <= _field_stack_stack_num_field_type_10_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h1 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_1_field_type_10_sub_class_id <= _field_stack_stack_num_field_type_10_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h1 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_1_field_type_11_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_11_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h1 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_1_field_type_11_field_type <= _field_stack_stack_num_field_type_11_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h1 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_1_field_type_11_sub_class_id <= _field_stack_stack_num_field_type_11_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h1 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_1_field_type_12_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_12_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h1 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_1_field_type_12_field_type <= _field_stack_stack_num_field_type_12_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h1 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_1_field_type_12_sub_class_id <= _field_stack_stack_num_field_type_12_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h1 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_1_field_type_13_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_13_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h1 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_1_field_type_13_field_type <= _field_stack_stack_num_field_type_13_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h1 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_1_field_type_13_sub_class_id <= _field_stack_stack_num_field_type_13_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h1 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_1_field_type_14_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_14_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h1 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_1_field_type_14_field_type <= _field_stack_stack_num_field_type_14_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h1 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_1_field_type_14_sub_class_id <= _field_stack_stack_num_field_type_14_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h1 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_1_field_type_15_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_15_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h1 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_1_field_type_15_field_type <= _field_stack_stack_num_field_type_15_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h1 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_1_field_type_15_sub_class_id <= _field_stack_stack_num_field_type_15_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h1 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_1_field_type_16_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_16_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h1 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_1_field_type_16_field_type <= _field_stack_stack_num_field_type_16_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h1 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_1_field_type_16_sub_class_id <= _field_stack_stack_num_field_type_16_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h1 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_1_field_type_17_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_17_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h1 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_1_field_type_17_field_type <= _field_stack_stack_num_field_type_17_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h1 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_1_field_type_17_sub_class_id <= _field_stack_stack_num_field_type_17_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h1 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_1_field_type_18_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_18_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h1 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_1_field_type_18_field_type <= _field_stack_stack_num_field_type_18_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h1 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_1_field_type_18_sub_class_id <= _field_stack_stack_num_field_type_18_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h1 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_1_field_type_19_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_19_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h1 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_1_field_type_19_field_type <= _field_stack_stack_num_field_type_19_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h1 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_1_field_type_19_sub_class_id <= _field_stack_stack_num_field_type_19_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h1 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_1_field_type_20_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_20_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h1 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_1_field_type_20_field_type <= _field_stack_stack_num_field_type_20_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h1 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_1_field_type_20_sub_class_id <= _field_stack_stack_num_field_type_20_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h1 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_1_field_type_21_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_21_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h1 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_1_field_type_21_field_type <= _field_stack_stack_num_field_type_21_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h1 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_1_field_type_21_sub_class_id <= _field_stack_stack_num_field_type_21_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h1 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_1_field_type_22_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_22_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h1 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_1_field_type_22_field_type <= _field_stack_stack_num_field_type_22_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h1 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_1_field_type_22_sub_class_id <= _field_stack_stack_num_field_type_22_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h1 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_1_field_type_23_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_23_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h1 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_1_field_type_23_field_type <= _field_stack_stack_num_field_type_23_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h1 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_1_field_type_23_sub_class_id <= _field_stack_stack_num_field_type_23_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h1 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_1_field_type_24_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_24_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h1 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_1_field_type_24_field_type <= _field_stack_stack_num_field_type_24_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h1 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_1_field_type_24_sub_class_id <= _field_stack_stack_num_field_type_24_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h1 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_1_field_type_25_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_25_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h1 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_1_field_type_25_field_type <= _field_stack_stack_num_field_type_25_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h1 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_1_field_type_25_sub_class_id <= _field_stack_stack_num_field_type_25_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h1 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_1_field_type_26_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_26_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h1 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_1_field_type_26_field_type <= _field_stack_stack_num_field_type_26_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h1 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_1_field_type_26_sub_class_id <= _field_stack_stack_num_field_type_26_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h1 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_1_field_type_27_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_27_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h1 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_1_field_type_27_field_type <= _field_stack_stack_num_field_type_27_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h1 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_1_field_type_27_sub_class_id <= _field_stack_stack_num_field_type_27_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h1 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_1_field_type_28_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_28_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h1 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_1_field_type_28_field_type <= _field_stack_stack_num_field_type_28_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h1 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_1_field_type_28_sub_class_id <= _field_stack_stack_num_field_type_28_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h1 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_1_field_type_29_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_29_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h1 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_1_field_type_29_field_type <= _field_stack_stack_num_field_type_29_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h1 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_1_field_type_29_sub_class_id <= _field_stack_stack_num_field_type_29_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h1 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_1_field_type_30_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_30_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h1 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_1_field_type_30_field_type <= _field_stack_stack_num_field_type_30_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h1 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_1_field_type_30_sub_class_id <= _field_stack_stack_num_field_type_30_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h1 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_1_field_type_31_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_31_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h1 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_1_field_type_31_field_type <= _field_stack_stack_num_field_type_31_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h1 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_1_field_type_31_sub_class_id <= _field_stack_stack_num_field_type_31_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h1 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_1_field_type_32_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_32_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h1 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_1_field_type_32_field_type <= _field_stack_stack_num_field_type_32_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h1 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_1_field_type_32_sub_class_id <= _field_stack_stack_num_field_type_32_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h2 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_2_field_type_0_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_0_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h2 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_2_field_type_0_field_type <= _field_stack_stack_num_field_type_0_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h2 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_2_field_type_0_sub_class_id <= _field_stack_stack_num_field_type_0_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h2 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_2_field_type_1_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_1_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h2 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_2_field_type_1_field_type <= _field_stack_stack_num_field_type_1_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h2 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_2_field_type_1_sub_class_id <= _field_stack_stack_num_field_type_1_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h2 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_2_field_type_2_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_2_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h2 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_2_field_type_2_field_type <= _field_stack_stack_num_field_type_2_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h2 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_2_field_type_2_sub_class_id <= _field_stack_stack_num_field_type_2_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h2 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_2_field_type_3_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_3_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h2 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_2_field_type_3_field_type <= _field_stack_stack_num_field_type_3_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h2 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_2_field_type_3_sub_class_id <= _field_stack_stack_num_field_type_3_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h2 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_2_field_type_4_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_4_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h2 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_2_field_type_4_field_type <= _field_stack_stack_num_field_type_4_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h2 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_2_field_type_4_sub_class_id <= _field_stack_stack_num_field_type_4_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h2 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_2_field_type_5_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_5_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h2 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_2_field_type_5_field_type <= _field_stack_stack_num_field_type_5_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h2 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_2_field_type_5_sub_class_id <= _field_stack_stack_num_field_type_5_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h2 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_2_field_type_6_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_6_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h2 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_2_field_type_6_field_type <= _field_stack_stack_num_field_type_6_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h2 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_2_field_type_6_sub_class_id <= _field_stack_stack_num_field_type_6_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h2 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_2_field_type_7_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_7_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h2 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_2_field_type_7_field_type <= _field_stack_stack_num_field_type_7_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h2 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_2_field_type_7_sub_class_id <= _field_stack_stack_num_field_type_7_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h2 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_2_field_type_8_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_8_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h2 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_2_field_type_8_field_type <= _field_stack_stack_num_field_type_8_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h2 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_2_field_type_8_sub_class_id <= _field_stack_stack_num_field_type_8_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h2 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_2_field_type_9_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_9_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h2 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_2_field_type_9_field_type <= _field_stack_stack_num_field_type_9_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h2 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_2_field_type_9_sub_class_id <= _field_stack_stack_num_field_type_9_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h2 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_2_field_type_10_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_10_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h2 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_2_field_type_10_field_type <= _field_stack_stack_num_field_type_10_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h2 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_2_field_type_10_sub_class_id <= _field_stack_stack_num_field_type_10_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h2 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_2_field_type_11_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_11_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h2 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_2_field_type_11_field_type <= _field_stack_stack_num_field_type_11_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h2 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_2_field_type_11_sub_class_id <= _field_stack_stack_num_field_type_11_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h2 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_2_field_type_12_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_12_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h2 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_2_field_type_12_field_type <= _field_stack_stack_num_field_type_12_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h2 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_2_field_type_12_sub_class_id <= _field_stack_stack_num_field_type_12_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h2 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_2_field_type_13_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_13_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h2 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_2_field_type_13_field_type <= _field_stack_stack_num_field_type_13_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h2 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_2_field_type_13_sub_class_id <= _field_stack_stack_num_field_type_13_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h2 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_2_field_type_14_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_14_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h2 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_2_field_type_14_field_type <= _field_stack_stack_num_field_type_14_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h2 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_2_field_type_14_sub_class_id <= _field_stack_stack_num_field_type_14_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h2 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_2_field_type_15_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_15_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h2 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_2_field_type_15_field_type <= _field_stack_stack_num_field_type_15_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h2 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_2_field_type_15_sub_class_id <= _field_stack_stack_num_field_type_15_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h2 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_2_field_type_16_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_16_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h2 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_2_field_type_16_field_type <= _field_stack_stack_num_field_type_16_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h2 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_2_field_type_16_sub_class_id <= _field_stack_stack_num_field_type_16_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h2 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_2_field_type_17_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_17_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h2 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_2_field_type_17_field_type <= _field_stack_stack_num_field_type_17_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h2 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_2_field_type_17_sub_class_id <= _field_stack_stack_num_field_type_17_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h2 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_2_field_type_18_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_18_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h2 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_2_field_type_18_field_type <= _field_stack_stack_num_field_type_18_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h2 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_2_field_type_18_sub_class_id <= _field_stack_stack_num_field_type_18_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h2 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_2_field_type_19_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_19_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h2 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_2_field_type_19_field_type <= _field_stack_stack_num_field_type_19_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h2 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_2_field_type_19_sub_class_id <= _field_stack_stack_num_field_type_19_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h2 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_2_field_type_20_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_20_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h2 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_2_field_type_20_field_type <= _field_stack_stack_num_field_type_20_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h2 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_2_field_type_20_sub_class_id <= _field_stack_stack_num_field_type_20_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h2 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_2_field_type_21_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_21_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h2 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_2_field_type_21_field_type <= _field_stack_stack_num_field_type_21_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h2 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_2_field_type_21_sub_class_id <= _field_stack_stack_num_field_type_21_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h2 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_2_field_type_22_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_22_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h2 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_2_field_type_22_field_type <= _field_stack_stack_num_field_type_22_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h2 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_2_field_type_22_sub_class_id <= _field_stack_stack_num_field_type_22_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h2 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_2_field_type_23_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_23_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h2 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_2_field_type_23_field_type <= _field_stack_stack_num_field_type_23_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h2 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_2_field_type_23_sub_class_id <= _field_stack_stack_num_field_type_23_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h2 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_2_field_type_24_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_24_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h2 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_2_field_type_24_field_type <= _field_stack_stack_num_field_type_24_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h2 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_2_field_type_24_sub_class_id <= _field_stack_stack_num_field_type_24_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h2 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_2_field_type_25_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_25_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h2 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_2_field_type_25_field_type <= _field_stack_stack_num_field_type_25_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h2 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_2_field_type_25_sub_class_id <= _field_stack_stack_num_field_type_25_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h2 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_2_field_type_26_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_26_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h2 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_2_field_type_26_field_type <= _field_stack_stack_num_field_type_26_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h2 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_2_field_type_26_sub_class_id <= _field_stack_stack_num_field_type_26_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h2 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_2_field_type_27_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_27_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h2 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_2_field_type_27_field_type <= _field_stack_stack_num_field_type_27_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h2 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_2_field_type_27_sub_class_id <= _field_stack_stack_num_field_type_27_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h2 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_2_field_type_28_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_28_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h2 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_2_field_type_28_field_type <= _field_stack_stack_num_field_type_28_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h2 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_2_field_type_28_sub_class_id <= _field_stack_stack_num_field_type_28_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h2 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_2_field_type_29_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_29_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h2 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_2_field_type_29_field_type <= _field_stack_stack_num_field_type_29_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h2 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_2_field_type_29_sub_class_id <= _field_stack_stack_num_field_type_29_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h2 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_2_field_type_30_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_30_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h2 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_2_field_type_30_field_type <= _field_stack_stack_num_field_type_30_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h2 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_2_field_type_30_sub_class_id <= _field_stack_stack_num_field_type_30_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h2 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_2_field_type_31_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_31_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h2 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_2_field_type_31_field_type <= _field_stack_stack_num_field_type_31_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h2 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_2_field_type_31_sub_class_id <= _field_stack_stack_num_field_type_31_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h2 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_2_field_type_32_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_32_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h2 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_2_field_type_32_field_type <= _field_stack_stack_num_field_type_32_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h2 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_2_field_type_32_sub_class_id <= _field_stack_stack_num_field_type_32_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h3 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_3_field_type_0_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_0_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h3 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_3_field_type_0_field_type <= _field_stack_stack_num_field_type_0_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h3 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_3_field_type_0_sub_class_id <= _field_stack_stack_num_field_type_0_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h3 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_3_field_type_1_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_1_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h3 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_3_field_type_1_field_type <= _field_stack_stack_num_field_type_1_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h3 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_3_field_type_1_sub_class_id <= _field_stack_stack_num_field_type_1_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h3 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_3_field_type_2_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_2_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h3 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_3_field_type_2_field_type <= _field_stack_stack_num_field_type_2_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h3 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_3_field_type_2_sub_class_id <= _field_stack_stack_num_field_type_2_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h3 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_3_field_type_3_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_3_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h3 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_3_field_type_3_field_type <= _field_stack_stack_num_field_type_3_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h3 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_3_field_type_3_sub_class_id <= _field_stack_stack_num_field_type_3_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h3 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_3_field_type_4_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_4_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h3 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_3_field_type_4_field_type <= _field_stack_stack_num_field_type_4_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h3 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_3_field_type_4_sub_class_id <= _field_stack_stack_num_field_type_4_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h3 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_3_field_type_5_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_5_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h3 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_3_field_type_5_field_type <= _field_stack_stack_num_field_type_5_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h3 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_3_field_type_5_sub_class_id <= _field_stack_stack_num_field_type_5_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h3 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_3_field_type_6_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_6_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h3 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_3_field_type_6_field_type <= _field_stack_stack_num_field_type_6_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h3 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_3_field_type_6_sub_class_id <= _field_stack_stack_num_field_type_6_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h3 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_3_field_type_7_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_7_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h3 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_3_field_type_7_field_type <= _field_stack_stack_num_field_type_7_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h3 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_3_field_type_7_sub_class_id <= _field_stack_stack_num_field_type_7_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h3 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_3_field_type_8_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_8_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h3 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_3_field_type_8_field_type <= _field_stack_stack_num_field_type_8_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h3 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_3_field_type_8_sub_class_id <= _field_stack_stack_num_field_type_8_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h3 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_3_field_type_9_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_9_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h3 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_3_field_type_9_field_type <= _field_stack_stack_num_field_type_9_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h3 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_3_field_type_9_sub_class_id <= _field_stack_stack_num_field_type_9_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h3 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_3_field_type_10_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_10_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h3 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_3_field_type_10_field_type <= _field_stack_stack_num_field_type_10_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h3 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_3_field_type_10_sub_class_id <= _field_stack_stack_num_field_type_10_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h3 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_3_field_type_11_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_11_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h3 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_3_field_type_11_field_type <= _field_stack_stack_num_field_type_11_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h3 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_3_field_type_11_sub_class_id <= _field_stack_stack_num_field_type_11_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h3 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_3_field_type_12_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_12_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h3 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_3_field_type_12_field_type <= _field_stack_stack_num_field_type_12_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h3 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_3_field_type_12_sub_class_id <= _field_stack_stack_num_field_type_12_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h3 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_3_field_type_13_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_13_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h3 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_3_field_type_13_field_type <= _field_stack_stack_num_field_type_13_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h3 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_3_field_type_13_sub_class_id <= _field_stack_stack_num_field_type_13_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h3 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_3_field_type_14_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_14_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h3 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_3_field_type_14_field_type <= _field_stack_stack_num_field_type_14_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h3 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_3_field_type_14_sub_class_id <= _field_stack_stack_num_field_type_14_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h3 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_3_field_type_15_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_15_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h3 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_3_field_type_15_field_type <= _field_stack_stack_num_field_type_15_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h3 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_3_field_type_15_sub_class_id <= _field_stack_stack_num_field_type_15_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h3 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_3_field_type_16_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_16_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h3 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_3_field_type_16_field_type <= _field_stack_stack_num_field_type_16_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h3 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_3_field_type_16_sub_class_id <= _field_stack_stack_num_field_type_16_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h3 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_3_field_type_17_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_17_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h3 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_3_field_type_17_field_type <= _field_stack_stack_num_field_type_17_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h3 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_3_field_type_17_sub_class_id <= _field_stack_stack_num_field_type_17_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h3 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_3_field_type_18_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_18_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h3 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_3_field_type_18_field_type <= _field_stack_stack_num_field_type_18_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h3 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_3_field_type_18_sub_class_id <= _field_stack_stack_num_field_type_18_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h3 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_3_field_type_19_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_19_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h3 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_3_field_type_19_field_type <= _field_stack_stack_num_field_type_19_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h3 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_3_field_type_19_sub_class_id <= _field_stack_stack_num_field_type_19_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h3 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_3_field_type_20_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_20_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h3 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_3_field_type_20_field_type <= _field_stack_stack_num_field_type_20_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h3 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_3_field_type_20_sub_class_id <= _field_stack_stack_num_field_type_20_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h3 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_3_field_type_21_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_21_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h3 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_3_field_type_21_field_type <= _field_stack_stack_num_field_type_21_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h3 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_3_field_type_21_sub_class_id <= _field_stack_stack_num_field_type_21_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h3 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_3_field_type_22_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_22_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h3 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_3_field_type_22_field_type <= _field_stack_stack_num_field_type_22_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h3 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_3_field_type_22_sub_class_id <= _field_stack_stack_num_field_type_22_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h3 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_3_field_type_23_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_23_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h3 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_3_field_type_23_field_type <= _field_stack_stack_num_field_type_23_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h3 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_3_field_type_23_sub_class_id <= _field_stack_stack_num_field_type_23_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h3 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_3_field_type_24_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_24_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h3 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_3_field_type_24_field_type <= _field_stack_stack_num_field_type_24_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h3 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_3_field_type_24_sub_class_id <= _field_stack_stack_num_field_type_24_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h3 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_3_field_type_25_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_25_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h3 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_3_field_type_25_field_type <= _field_stack_stack_num_field_type_25_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h3 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_3_field_type_25_sub_class_id <= _field_stack_stack_num_field_type_25_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h3 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_3_field_type_26_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_26_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h3 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_3_field_type_26_field_type <= _field_stack_stack_num_field_type_26_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h3 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_3_field_type_26_sub_class_id <= _field_stack_stack_num_field_type_26_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h3 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_3_field_type_27_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_27_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h3 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_3_field_type_27_field_type <= _field_stack_stack_num_field_type_27_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h3 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_3_field_type_27_sub_class_id <= _field_stack_stack_num_field_type_27_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h3 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_3_field_type_28_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_28_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h3 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_3_field_type_28_field_type <= _field_stack_stack_num_field_type_28_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h3 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_3_field_type_28_sub_class_id <= _field_stack_stack_num_field_type_28_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h3 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_3_field_type_29_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_29_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h3 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_3_field_type_29_field_type <= _field_stack_stack_num_field_type_29_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h3 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_3_field_type_29_sub_class_id <= _field_stack_stack_num_field_type_29_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h3 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_3_field_type_30_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_30_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h3 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_3_field_type_30_field_type <= _field_stack_stack_num_field_type_30_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h3 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_3_field_type_30_sub_class_id <= _field_stack_stack_num_field_type_30_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h3 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_3_field_type_31_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_31_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h3 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_3_field_type_31_field_type <= _field_stack_stack_num_field_type_31_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h3 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_3_field_type_31_sub_class_id <= _field_stack_stack_num_field_type_31_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h3 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_3_field_type_32_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_32_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h3 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_3_field_type_32_field_type <= _field_stack_stack_num_field_type_32_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h3 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_3_field_type_32_sub_class_id <= _field_stack_stack_num_field_type_32_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h4 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_4_field_type_0_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_0_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h4 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_4_field_type_0_field_type <= _field_stack_stack_num_field_type_0_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h4 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_4_field_type_0_sub_class_id <= _field_stack_stack_num_field_type_0_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h4 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_4_field_type_1_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_1_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h4 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_4_field_type_1_field_type <= _field_stack_stack_num_field_type_1_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h4 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_4_field_type_1_sub_class_id <= _field_stack_stack_num_field_type_1_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h4 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_4_field_type_2_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_2_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h4 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_4_field_type_2_field_type <= _field_stack_stack_num_field_type_2_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h4 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_4_field_type_2_sub_class_id <= _field_stack_stack_num_field_type_2_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h4 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_4_field_type_3_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_3_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h4 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_4_field_type_3_field_type <= _field_stack_stack_num_field_type_3_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h4 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_4_field_type_3_sub_class_id <= _field_stack_stack_num_field_type_3_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h4 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_4_field_type_4_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_4_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h4 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_4_field_type_4_field_type <= _field_stack_stack_num_field_type_4_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h4 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_4_field_type_4_sub_class_id <= _field_stack_stack_num_field_type_4_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h4 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_4_field_type_5_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_5_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h4 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_4_field_type_5_field_type <= _field_stack_stack_num_field_type_5_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h4 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_4_field_type_5_sub_class_id <= _field_stack_stack_num_field_type_5_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h4 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_4_field_type_6_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_6_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h4 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_4_field_type_6_field_type <= _field_stack_stack_num_field_type_6_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h4 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_4_field_type_6_sub_class_id <= _field_stack_stack_num_field_type_6_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h4 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_4_field_type_7_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_7_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h4 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_4_field_type_7_field_type <= _field_stack_stack_num_field_type_7_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h4 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_4_field_type_7_sub_class_id <= _field_stack_stack_num_field_type_7_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h4 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_4_field_type_8_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_8_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h4 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_4_field_type_8_field_type <= _field_stack_stack_num_field_type_8_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h4 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_4_field_type_8_sub_class_id <= _field_stack_stack_num_field_type_8_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h4 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_4_field_type_9_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_9_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h4 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_4_field_type_9_field_type <= _field_stack_stack_num_field_type_9_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h4 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_4_field_type_9_sub_class_id <= _field_stack_stack_num_field_type_9_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h4 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_4_field_type_10_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_10_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h4 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_4_field_type_10_field_type <= _field_stack_stack_num_field_type_10_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h4 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_4_field_type_10_sub_class_id <= _field_stack_stack_num_field_type_10_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h4 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_4_field_type_11_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_11_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h4 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_4_field_type_11_field_type <= _field_stack_stack_num_field_type_11_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h4 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_4_field_type_11_sub_class_id <= _field_stack_stack_num_field_type_11_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h4 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_4_field_type_12_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_12_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h4 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_4_field_type_12_field_type <= _field_stack_stack_num_field_type_12_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h4 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_4_field_type_12_sub_class_id <= _field_stack_stack_num_field_type_12_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h4 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_4_field_type_13_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_13_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h4 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_4_field_type_13_field_type <= _field_stack_stack_num_field_type_13_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h4 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_4_field_type_13_sub_class_id <= _field_stack_stack_num_field_type_13_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h4 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_4_field_type_14_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_14_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h4 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_4_field_type_14_field_type <= _field_stack_stack_num_field_type_14_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h4 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_4_field_type_14_sub_class_id <= _field_stack_stack_num_field_type_14_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h4 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_4_field_type_15_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_15_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h4 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_4_field_type_15_field_type <= _field_stack_stack_num_field_type_15_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h4 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_4_field_type_15_sub_class_id <= _field_stack_stack_num_field_type_15_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h4 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_4_field_type_16_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_16_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h4 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_4_field_type_16_field_type <= _field_stack_stack_num_field_type_16_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h4 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_4_field_type_16_sub_class_id <= _field_stack_stack_num_field_type_16_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h4 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_4_field_type_17_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_17_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h4 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_4_field_type_17_field_type <= _field_stack_stack_num_field_type_17_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h4 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_4_field_type_17_sub_class_id <= _field_stack_stack_num_field_type_17_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h4 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_4_field_type_18_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_18_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h4 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_4_field_type_18_field_type <= _field_stack_stack_num_field_type_18_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h4 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_4_field_type_18_sub_class_id <= _field_stack_stack_num_field_type_18_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h4 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_4_field_type_19_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_19_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h4 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_4_field_type_19_field_type <= _field_stack_stack_num_field_type_19_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h4 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_4_field_type_19_sub_class_id <= _field_stack_stack_num_field_type_19_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h4 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_4_field_type_20_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_20_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h4 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_4_field_type_20_field_type <= _field_stack_stack_num_field_type_20_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h4 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_4_field_type_20_sub_class_id <= _field_stack_stack_num_field_type_20_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h4 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_4_field_type_21_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_21_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h4 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_4_field_type_21_field_type <= _field_stack_stack_num_field_type_21_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h4 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_4_field_type_21_sub_class_id <= _field_stack_stack_num_field_type_21_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h4 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_4_field_type_22_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_22_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h4 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_4_field_type_22_field_type <= _field_stack_stack_num_field_type_22_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h4 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_4_field_type_22_sub_class_id <= _field_stack_stack_num_field_type_22_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h4 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_4_field_type_23_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_23_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h4 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_4_field_type_23_field_type <= _field_stack_stack_num_field_type_23_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h4 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_4_field_type_23_sub_class_id <= _field_stack_stack_num_field_type_23_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h4 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_4_field_type_24_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_24_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h4 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_4_field_type_24_field_type <= _field_stack_stack_num_field_type_24_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h4 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_4_field_type_24_sub_class_id <= _field_stack_stack_num_field_type_24_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h4 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_4_field_type_25_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_25_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h4 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_4_field_type_25_field_type <= _field_stack_stack_num_field_type_25_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h4 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_4_field_type_25_sub_class_id <= _field_stack_stack_num_field_type_25_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h4 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_4_field_type_26_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_26_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h4 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_4_field_type_26_field_type <= _field_stack_stack_num_field_type_26_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h4 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_4_field_type_26_sub_class_id <= _field_stack_stack_num_field_type_26_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h4 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_4_field_type_27_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_27_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h4 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_4_field_type_27_field_type <= _field_stack_stack_num_field_type_27_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h4 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_4_field_type_27_sub_class_id <= _field_stack_stack_num_field_type_27_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h4 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_4_field_type_28_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_28_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h4 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_4_field_type_28_field_type <= _field_stack_stack_num_field_type_28_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h4 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_4_field_type_28_sub_class_id <= _field_stack_stack_num_field_type_28_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h4 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_4_field_type_29_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_29_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h4 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_4_field_type_29_field_type <= _field_stack_stack_num_field_type_29_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h4 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_4_field_type_29_sub_class_id <= _field_stack_stack_num_field_type_29_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h4 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_4_field_type_30_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_30_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h4 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_4_field_type_30_field_type <= _field_stack_stack_num_field_type_30_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h4 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_4_field_type_30_sub_class_id <= _field_stack_stack_num_field_type_30_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h4 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_4_field_type_31_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_31_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h4 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_4_field_type_31_field_type <= _field_stack_stack_num_field_type_31_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h4 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_4_field_type_31_sub_class_id <= _field_stack_stack_num_field_type_31_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h4 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_4_field_type_32_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_32_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h4 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_4_field_type_32_field_type <= _field_stack_stack_num_field_type_32_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h4 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_4_field_type_32_sub_class_id <= _field_stack_stack_num_field_type_32_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h5 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_5_field_type_0_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_0_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h5 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_5_field_type_0_field_type <= _field_stack_stack_num_field_type_0_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h5 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_5_field_type_0_sub_class_id <= _field_stack_stack_num_field_type_0_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h5 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_5_field_type_1_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_1_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h5 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_5_field_type_1_field_type <= _field_stack_stack_num_field_type_1_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h5 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_5_field_type_1_sub_class_id <= _field_stack_stack_num_field_type_1_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h5 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_5_field_type_2_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_2_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h5 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_5_field_type_2_field_type <= _field_stack_stack_num_field_type_2_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h5 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_5_field_type_2_sub_class_id <= _field_stack_stack_num_field_type_2_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h5 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_5_field_type_3_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_3_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h5 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_5_field_type_3_field_type <= _field_stack_stack_num_field_type_3_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h5 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_5_field_type_3_sub_class_id <= _field_stack_stack_num_field_type_3_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h5 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_5_field_type_4_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_4_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h5 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_5_field_type_4_field_type <= _field_stack_stack_num_field_type_4_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h5 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_5_field_type_4_sub_class_id <= _field_stack_stack_num_field_type_4_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h5 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_5_field_type_5_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_5_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h5 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_5_field_type_5_field_type <= _field_stack_stack_num_field_type_5_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h5 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_5_field_type_5_sub_class_id <= _field_stack_stack_num_field_type_5_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h5 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_5_field_type_6_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_6_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h5 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_5_field_type_6_field_type <= _field_stack_stack_num_field_type_6_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h5 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_5_field_type_6_sub_class_id <= _field_stack_stack_num_field_type_6_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h5 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_5_field_type_7_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_7_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h5 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_5_field_type_7_field_type <= _field_stack_stack_num_field_type_7_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h5 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_5_field_type_7_sub_class_id <= _field_stack_stack_num_field_type_7_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h5 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_5_field_type_8_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_8_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h5 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_5_field_type_8_field_type <= _field_stack_stack_num_field_type_8_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h5 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_5_field_type_8_sub_class_id <= _field_stack_stack_num_field_type_8_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h5 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_5_field_type_9_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_9_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h5 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_5_field_type_9_field_type <= _field_stack_stack_num_field_type_9_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h5 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_5_field_type_9_sub_class_id <= _field_stack_stack_num_field_type_9_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h5 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_5_field_type_10_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_10_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h5 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_5_field_type_10_field_type <= _field_stack_stack_num_field_type_10_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h5 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_5_field_type_10_sub_class_id <= _field_stack_stack_num_field_type_10_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h5 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_5_field_type_11_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_11_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h5 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_5_field_type_11_field_type <= _field_stack_stack_num_field_type_11_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h5 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_5_field_type_11_sub_class_id <= _field_stack_stack_num_field_type_11_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h5 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_5_field_type_12_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_12_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h5 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_5_field_type_12_field_type <= _field_stack_stack_num_field_type_12_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h5 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_5_field_type_12_sub_class_id <= _field_stack_stack_num_field_type_12_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h5 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_5_field_type_13_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_13_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h5 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_5_field_type_13_field_type <= _field_stack_stack_num_field_type_13_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h5 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_5_field_type_13_sub_class_id <= _field_stack_stack_num_field_type_13_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h5 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_5_field_type_14_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_14_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h5 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_5_field_type_14_field_type <= _field_stack_stack_num_field_type_14_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h5 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_5_field_type_14_sub_class_id <= _field_stack_stack_num_field_type_14_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h5 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_5_field_type_15_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_15_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h5 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_5_field_type_15_field_type <= _field_stack_stack_num_field_type_15_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h5 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_5_field_type_15_sub_class_id <= _field_stack_stack_num_field_type_15_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h5 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_5_field_type_16_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_16_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h5 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_5_field_type_16_field_type <= _field_stack_stack_num_field_type_16_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h5 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_5_field_type_16_sub_class_id <= _field_stack_stack_num_field_type_16_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h5 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_5_field_type_17_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_17_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h5 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_5_field_type_17_field_type <= _field_stack_stack_num_field_type_17_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h5 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_5_field_type_17_sub_class_id <= _field_stack_stack_num_field_type_17_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h5 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_5_field_type_18_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_18_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h5 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_5_field_type_18_field_type <= _field_stack_stack_num_field_type_18_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h5 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_5_field_type_18_sub_class_id <= _field_stack_stack_num_field_type_18_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h5 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_5_field_type_19_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_19_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h5 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_5_field_type_19_field_type <= _field_stack_stack_num_field_type_19_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h5 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_5_field_type_19_sub_class_id <= _field_stack_stack_num_field_type_19_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h5 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_5_field_type_20_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_20_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h5 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_5_field_type_20_field_type <= _field_stack_stack_num_field_type_20_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h5 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_5_field_type_20_sub_class_id <= _field_stack_stack_num_field_type_20_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h5 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_5_field_type_21_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_21_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h5 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_5_field_type_21_field_type <= _field_stack_stack_num_field_type_21_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h5 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_5_field_type_21_sub_class_id <= _field_stack_stack_num_field_type_21_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h5 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_5_field_type_22_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_22_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h5 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_5_field_type_22_field_type <= _field_stack_stack_num_field_type_22_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h5 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_5_field_type_22_sub_class_id <= _field_stack_stack_num_field_type_22_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h5 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_5_field_type_23_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_23_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h5 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_5_field_type_23_field_type <= _field_stack_stack_num_field_type_23_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h5 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_5_field_type_23_sub_class_id <= _field_stack_stack_num_field_type_23_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h5 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_5_field_type_24_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_24_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h5 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_5_field_type_24_field_type <= _field_stack_stack_num_field_type_24_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h5 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_5_field_type_24_sub_class_id <= _field_stack_stack_num_field_type_24_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h5 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_5_field_type_25_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_25_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h5 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_5_field_type_25_field_type <= _field_stack_stack_num_field_type_25_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h5 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_5_field_type_25_sub_class_id <= _field_stack_stack_num_field_type_25_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h5 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_5_field_type_26_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_26_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h5 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_5_field_type_26_field_type <= _field_stack_stack_num_field_type_26_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h5 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_5_field_type_26_sub_class_id <= _field_stack_stack_num_field_type_26_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h5 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_5_field_type_27_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_27_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h5 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_5_field_type_27_field_type <= _field_stack_stack_num_field_type_27_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h5 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_5_field_type_27_sub_class_id <= _field_stack_stack_num_field_type_27_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h5 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_5_field_type_28_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_28_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h5 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_5_field_type_28_field_type <= _field_stack_stack_num_field_type_28_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h5 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_5_field_type_28_sub_class_id <= _field_stack_stack_num_field_type_28_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h5 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_5_field_type_29_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_29_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h5 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_5_field_type_29_field_type <= _field_stack_stack_num_field_type_29_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h5 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_5_field_type_29_sub_class_id <= _field_stack_stack_num_field_type_29_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h5 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_5_field_type_30_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_30_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h5 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_5_field_type_30_field_type <= _field_stack_stack_num_field_type_30_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h5 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_5_field_type_30_sub_class_id <= _field_stack_stack_num_field_type_30_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h5 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_5_field_type_31_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_31_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h5 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_5_field_type_31_field_type <= _field_stack_stack_num_field_type_31_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h5 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_5_field_type_31_sub_class_id <= _field_stack_stack_num_field_type_31_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h5 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_5_field_type_32_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_32_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h5 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_5_field_type_32_field_type <= _field_stack_stack_num_field_type_32_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h5 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_5_field_type_32_sub_class_id <= _field_stack_stack_num_field_type_32_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h6 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_6_field_type_0_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_0_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h6 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_6_field_type_0_field_type <= _field_stack_stack_num_field_type_0_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h6 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_6_field_type_0_sub_class_id <= _field_stack_stack_num_field_type_0_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h6 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_6_field_type_1_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_1_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h6 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_6_field_type_1_field_type <= _field_stack_stack_num_field_type_1_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h6 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_6_field_type_1_sub_class_id <= _field_stack_stack_num_field_type_1_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h6 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_6_field_type_2_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_2_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h6 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_6_field_type_2_field_type <= _field_stack_stack_num_field_type_2_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h6 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_6_field_type_2_sub_class_id <= _field_stack_stack_num_field_type_2_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h6 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_6_field_type_3_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_3_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h6 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_6_field_type_3_field_type <= _field_stack_stack_num_field_type_3_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h6 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_6_field_type_3_sub_class_id <= _field_stack_stack_num_field_type_3_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h6 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_6_field_type_4_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_4_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h6 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_6_field_type_4_field_type <= _field_stack_stack_num_field_type_4_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h6 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_6_field_type_4_sub_class_id <= _field_stack_stack_num_field_type_4_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h6 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_6_field_type_5_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_5_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h6 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_6_field_type_5_field_type <= _field_stack_stack_num_field_type_5_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h6 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_6_field_type_5_sub_class_id <= _field_stack_stack_num_field_type_5_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h6 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_6_field_type_6_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_6_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h6 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_6_field_type_6_field_type <= _field_stack_stack_num_field_type_6_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h6 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_6_field_type_6_sub_class_id <= _field_stack_stack_num_field_type_6_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h6 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_6_field_type_7_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_7_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h6 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_6_field_type_7_field_type <= _field_stack_stack_num_field_type_7_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h6 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_6_field_type_7_sub_class_id <= _field_stack_stack_num_field_type_7_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h6 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_6_field_type_8_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_8_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h6 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_6_field_type_8_field_type <= _field_stack_stack_num_field_type_8_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h6 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_6_field_type_8_sub_class_id <= _field_stack_stack_num_field_type_8_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h6 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_6_field_type_9_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_9_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h6 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_6_field_type_9_field_type <= _field_stack_stack_num_field_type_9_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h6 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_6_field_type_9_sub_class_id <= _field_stack_stack_num_field_type_9_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h6 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_6_field_type_10_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_10_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h6 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_6_field_type_10_field_type <= _field_stack_stack_num_field_type_10_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h6 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_6_field_type_10_sub_class_id <= _field_stack_stack_num_field_type_10_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h6 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_6_field_type_11_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_11_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h6 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_6_field_type_11_field_type <= _field_stack_stack_num_field_type_11_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h6 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_6_field_type_11_sub_class_id <= _field_stack_stack_num_field_type_11_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h6 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_6_field_type_12_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_12_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h6 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_6_field_type_12_field_type <= _field_stack_stack_num_field_type_12_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h6 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_6_field_type_12_sub_class_id <= _field_stack_stack_num_field_type_12_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h6 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_6_field_type_13_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_13_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h6 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_6_field_type_13_field_type <= _field_stack_stack_num_field_type_13_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h6 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_6_field_type_13_sub_class_id <= _field_stack_stack_num_field_type_13_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h6 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_6_field_type_14_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_14_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h6 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_6_field_type_14_field_type <= _field_stack_stack_num_field_type_14_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h6 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_6_field_type_14_sub_class_id <= _field_stack_stack_num_field_type_14_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h6 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_6_field_type_15_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_15_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h6 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_6_field_type_15_field_type <= _field_stack_stack_num_field_type_15_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h6 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_6_field_type_15_sub_class_id <= _field_stack_stack_num_field_type_15_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h6 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_6_field_type_16_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_16_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h6 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_6_field_type_16_field_type <= _field_stack_stack_num_field_type_16_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h6 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_6_field_type_16_sub_class_id <= _field_stack_stack_num_field_type_16_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h6 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_6_field_type_17_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_17_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h6 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_6_field_type_17_field_type <= _field_stack_stack_num_field_type_17_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h6 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_6_field_type_17_sub_class_id <= _field_stack_stack_num_field_type_17_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h6 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_6_field_type_18_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_18_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h6 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_6_field_type_18_field_type <= _field_stack_stack_num_field_type_18_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h6 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_6_field_type_18_sub_class_id <= _field_stack_stack_num_field_type_18_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h6 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_6_field_type_19_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_19_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h6 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_6_field_type_19_field_type <= _field_stack_stack_num_field_type_19_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h6 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_6_field_type_19_sub_class_id <= _field_stack_stack_num_field_type_19_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h6 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_6_field_type_20_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_20_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h6 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_6_field_type_20_field_type <= _field_stack_stack_num_field_type_20_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h6 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_6_field_type_20_sub_class_id <= _field_stack_stack_num_field_type_20_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h6 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_6_field_type_21_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_21_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h6 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_6_field_type_21_field_type <= _field_stack_stack_num_field_type_21_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h6 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_6_field_type_21_sub_class_id <= _field_stack_stack_num_field_type_21_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h6 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_6_field_type_22_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_22_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h6 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_6_field_type_22_field_type <= _field_stack_stack_num_field_type_22_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h6 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_6_field_type_22_sub_class_id <= _field_stack_stack_num_field_type_22_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h6 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_6_field_type_23_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_23_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h6 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_6_field_type_23_field_type <= _field_stack_stack_num_field_type_23_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h6 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_6_field_type_23_sub_class_id <= _field_stack_stack_num_field_type_23_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h6 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_6_field_type_24_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_24_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h6 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_6_field_type_24_field_type <= _field_stack_stack_num_field_type_24_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h6 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_6_field_type_24_sub_class_id <= _field_stack_stack_num_field_type_24_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h6 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_6_field_type_25_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_25_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h6 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_6_field_type_25_field_type <= _field_stack_stack_num_field_type_25_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h6 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_6_field_type_25_sub_class_id <= _field_stack_stack_num_field_type_25_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h6 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_6_field_type_26_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_26_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h6 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_6_field_type_26_field_type <= _field_stack_stack_num_field_type_26_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h6 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_6_field_type_26_sub_class_id <= _field_stack_stack_num_field_type_26_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h6 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_6_field_type_27_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_27_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h6 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_6_field_type_27_field_type <= _field_stack_stack_num_field_type_27_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h6 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_6_field_type_27_sub_class_id <= _field_stack_stack_num_field_type_27_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h6 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_6_field_type_28_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_28_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h6 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_6_field_type_28_field_type <= _field_stack_stack_num_field_type_28_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h6 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_6_field_type_28_sub_class_id <= _field_stack_stack_num_field_type_28_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h6 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_6_field_type_29_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_29_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h6 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_6_field_type_29_field_type <= _field_stack_stack_num_field_type_29_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h6 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_6_field_type_29_sub_class_id <= _field_stack_stack_num_field_type_29_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h6 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_6_field_type_30_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_30_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h6 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_6_field_type_30_field_type <= _field_stack_stack_num_field_type_30_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h6 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_6_field_type_30_sub_class_id <= _field_stack_stack_num_field_type_30_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h6 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_6_field_type_31_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_31_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h6 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_6_field_type_31_field_type <= _field_stack_stack_num_field_type_31_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h6 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_6_field_type_31_sub_class_id <= _field_stack_stack_num_field_type_31_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h6 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_6_field_type_32_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_32_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h6 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_6_field_type_32_field_type <= _field_stack_stack_num_field_type_32_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h6 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_6_field_type_32_sub_class_id <= _field_stack_stack_num_field_type_32_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h7 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_7_field_type_0_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_0_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h7 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_7_field_type_0_field_type <= _field_stack_stack_num_field_type_0_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h7 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_7_field_type_0_sub_class_id <= _field_stack_stack_num_field_type_0_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h7 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_7_field_type_1_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_1_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h7 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_7_field_type_1_field_type <= _field_stack_stack_num_field_type_1_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h7 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_7_field_type_1_sub_class_id <= _field_stack_stack_num_field_type_1_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h7 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_7_field_type_2_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_2_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h7 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_7_field_type_2_field_type <= _field_stack_stack_num_field_type_2_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h7 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_7_field_type_2_sub_class_id <= _field_stack_stack_num_field_type_2_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h7 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_7_field_type_3_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_3_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h7 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_7_field_type_3_field_type <= _field_stack_stack_num_field_type_3_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h7 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_7_field_type_3_sub_class_id <= _field_stack_stack_num_field_type_3_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h7 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_7_field_type_4_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_4_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h7 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_7_field_type_4_field_type <= _field_stack_stack_num_field_type_4_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h7 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_7_field_type_4_sub_class_id <= _field_stack_stack_num_field_type_4_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h7 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_7_field_type_5_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_5_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h7 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_7_field_type_5_field_type <= _field_stack_stack_num_field_type_5_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h7 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_7_field_type_5_sub_class_id <= _field_stack_stack_num_field_type_5_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h7 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_7_field_type_6_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_6_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h7 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_7_field_type_6_field_type <= _field_stack_stack_num_field_type_6_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h7 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_7_field_type_6_sub_class_id <= _field_stack_stack_num_field_type_6_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h7 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_7_field_type_7_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_7_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h7 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_7_field_type_7_field_type <= _field_stack_stack_num_field_type_7_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h7 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_7_field_type_7_sub_class_id <= _field_stack_stack_num_field_type_7_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h7 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_7_field_type_8_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_8_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h7 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_7_field_type_8_field_type <= _field_stack_stack_num_field_type_8_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h7 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_7_field_type_8_sub_class_id <= _field_stack_stack_num_field_type_8_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h7 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_7_field_type_9_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_9_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h7 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_7_field_type_9_field_type <= _field_stack_stack_num_field_type_9_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h7 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_7_field_type_9_sub_class_id <= _field_stack_stack_num_field_type_9_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h7 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_7_field_type_10_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_10_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h7 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_7_field_type_10_field_type <= _field_stack_stack_num_field_type_10_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h7 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_7_field_type_10_sub_class_id <= _field_stack_stack_num_field_type_10_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h7 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_7_field_type_11_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_11_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h7 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_7_field_type_11_field_type <= _field_stack_stack_num_field_type_11_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h7 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_7_field_type_11_sub_class_id <= _field_stack_stack_num_field_type_11_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h7 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_7_field_type_12_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_12_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h7 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_7_field_type_12_field_type <= _field_stack_stack_num_field_type_12_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h7 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_7_field_type_12_sub_class_id <= _field_stack_stack_num_field_type_12_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h7 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_7_field_type_13_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_13_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h7 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_7_field_type_13_field_type <= _field_stack_stack_num_field_type_13_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h7 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_7_field_type_13_sub_class_id <= _field_stack_stack_num_field_type_13_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h7 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_7_field_type_14_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_14_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h7 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_7_field_type_14_field_type <= _field_stack_stack_num_field_type_14_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h7 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_7_field_type_14_sub_class_id <= _field_stack_stack_num_field_type_14_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h7 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_7_field_type_15_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_15_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h7 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_7_field_type_15_field_type <= _field_stack_stack_num_field_type_15_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h7 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_7_field_type_15_sub_class_id <= _field_stack_stack_num_field_type_15_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h7 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_7_field_type_16_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_16_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h7 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_7_field_type_16_field_type <= _field_stack_stack_num_field_type_16_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h7 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_7_field_type_16_sub_class_id <= _field_stack_stack_num_field_type_16_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h7 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_7_field_type_17_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_17_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h7 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_7_field_type_17_field_type <= _field_stack_stack_num_field_type_17_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h7 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_7_field_type_17_sub_class_id <= _field_stack_stack_num_field_type_17_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h7 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_7_field_type_18_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_18_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h7 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_7_field_type_18_field_type <= _field_stack_stack_num_field_type_18_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h7 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_7_field_type_18_sub_class_id <= _field_stack_stack_num_field_type_18_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h7 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_7_field_type_19_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_19_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h7 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_7_field_type_19_field_type <= _field_stack_stack_num_field_type_19_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h7 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_7_field_type_19_sub_class_id <= _field_stack_stack_num_field_type_19_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h7 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_7_field_type_20_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_20_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h7 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_7_field_type_20_field_type <= _field_stack_stack_num_field_type_20_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h7 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_7_field_type_20_sub_class_id <= _field_stack_stack_num_field_type_20_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h7 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_7_field_type_21_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_21_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h7 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_7_field_type_21_field_type <= _field_stack_stack_num_field_type_21_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h7 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_7_field_type_21_sub_class_id <= _field_stack_stack_num_field_type_21_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h7 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_7_field_type_22_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_22_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h7 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_7_field_type_22_field_type <= _field_stack_stack_num_field_type_22_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h7 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_7_field_type_22_sub_class_id <= _field_stack_stack_num_field_type_22_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h7 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_7_field_type_23_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_23_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h7 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_7_field_type_23_field_type <= _field_stack_stack_num_field_type_23_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h7 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_7_field_type_23_sub_class_id <= _field_stack_stack_num_field_type_23_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h7 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_7_field_type_24_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_24_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h7 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_7_field_type_24_field_type <= _field_stack_stack_num_field_type_24_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h7 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_7_field_type_24_sub_class_id <= _field_stack_stack_num_field_type_24_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h7 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_7_field_type_25_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_25_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h7 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_7_field_type_25_field_type <= _field_stack_stack_num_field_type_25_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h7 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_7_field_type_25_sub_class_id <= _field_stack_stack_num_field_type_25_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h7 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_7_field_type_26_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_26_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h7 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_7_field_type_26_field_type <= _field_stack_stack_num_field_type_26_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h7 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_7_field_type_26_sub_class_id <= _field_stack_stack_num_field_type_26_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h7 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_7_field_type_27_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_27_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h7 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_7_field_type_27_field_type <= _field_stack_stack_num_field_type_27_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h7 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_7_field_type_27_sub_class_id <= _field_stack_stack_num_field_type_27_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h7 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_7_field_type_28_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_28_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h7 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_7_field_type_28_field_type <= _field_stack_stack_num_field_type_28_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h7 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_7_field_type_28_sub_class_id <= _field_stack_stack_num_field_type_28_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h7 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_7_field_type_29_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_29_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h7 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_7_field_type_29_field_type <= _field_stack_stack_num_field_type_29_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h7 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_7_field_type_29_sub_class_id <= _field_stack_stack_num_field_type_29_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h7 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_7_field_type_30_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_30_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h7 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_7_field_type_30_field_type <= _field_stack_stack_num_field_type_30_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h7 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_7_field_type_30_sub_class_id <= _field_stack_stack_num_field_type_30_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h7 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_7_field_type_31_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_31_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h7 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_7_field_type_31_field_type <= _field_stack_stack_num_field_type_31_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h7 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_7_field_type_31_sub_class_id <= _field_stack_stack_num_field_type_31_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h7 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_7_field_type_32_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_32_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h7 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_7_field_type_32_field_type <= _field_stack_stack_num_field_type_32_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h7 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_7_field_type_32_sub_class_id <= _field_stack_stack_num_field_type_32_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h8 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_8_field_type_0_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_0_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h8 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_8_field_type_0_field_type <= _field_stack_stack_num_field_type_0_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h8 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_8_field_type_0_sub_class_id <= _field_stack_stack_num_field_type_0_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h8 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_8_field_type_1_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_1_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h8 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_8_field_type_1_field_type <= _field_stack_stack_num_field_type_1_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h8 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_8_field_type_1_sub_class_id <= _field_stack_stack_num_field_type_1_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h8 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_8_field_type_2_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_2_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h8 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_8_field_type_2_field_type <= _field_stack_stack_num_field_type_2_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h8 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_8_field_type_2_sub_class_id <= _field_stack_stack_num_field_type_2_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h8 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_8_field_type_3_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_3_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h8 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_8_field_type_3_field_type <= _field_stack_stack_num_field_type_3_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h8 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_8_field_type_3_sub_class_id <= _field_stack_stack_num_field_type_3_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h8 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_8_field_type_4_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_4_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h8 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_8_field_type_4_field_type <= _field_stack_stack_num_field_type_4_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h8 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_8_field_type_4_sub_class_id <= _field_stack_stack_num_field_type_4_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h8 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_8_field_type_5_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_5_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h8 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_8_field_type_5_field_type <= _field_stack_stack_num_field_type_5_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h8 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_8_field_type_5_sub_class_id <= _field_stack_stack_num_field_type_5_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h8 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_8_field_type_6_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_6_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h8 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_8_field_type_6_field_type <= _field_stack_stack_num_field_type_6_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h8 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_8_field_type_6_sub_class_id <= _field_stack_stack_num_field_type_6_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h8 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_8_field_type_7_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_7_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h8 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_8_field_type_7_field_type <= _field_stack_stack_num_field_type_7_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h8 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_8_field_type_7_sub_class_id <= _field_stack_stack_num_field_type_7_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h8 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_8_field_type_8_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_8_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h8 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_8_field_type_8_field_type <= _field_stack_stack_num_field_type_8_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h8 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_8_field_type_8_sub_class_id <= _field_stack_stack_num_field_type_8_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h8 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_8_field_type_9_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_9_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h8 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_8_field_type_9_field_type <= _field_stack_stack_num_field_type_9_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h8 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_8_field_type_9_sub_class_id <= _field_stack_stack_num_field_type_9_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h8 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_8_field_type_10_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_10_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h8 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_8_field_type_10_field_type <= _field_stack_stack_num_field_type_10_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h8 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_8_field_type_10_sub_class_id <= _field_stack_stack_num_field_type_10_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h8 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_8_field_type_11_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_11_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h8 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_8_field_type_11_field_type <= _field_stack_stack_num_field_type_11_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h8 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_8_field_type_11_sub_class_id <= _field_stack_stack_num_field_type_11_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h8 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_8_field_type_12_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_12_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h8 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_8_field_type_12_field_type <= _field_stack_stack_num_field_type_12_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h8 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_8_field_type_12_sub_class_id <= _field_stack_stack_num_field_type_12_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h8 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_8_field_type_13_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_13_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h8 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_8_field_type_13_field_type <= _field_stack_stack_num_field_type_13_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h8 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_8_field_type_13_sub_class_id <= _field_stack_stack_num_field_type_13_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h8 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_8_field_type_14_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_14_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h8 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_8_field_type_14_field_type <= _field_stack_stack_num_field_type_14_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h8 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_8_field_type_14_sub_class_id <= _field_stack_stack_num_field_type_14_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h8 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_8_field_type_15_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_15_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h8 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_8_field_type_15_field_type <= _field_stack_stack_num_field_type_15_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h8 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_8_field_type_15_sub_class_id <= _field_stack_stack_num_field_type_15_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h8 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_8_field_type_16_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_16_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h8 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_8_field_type_16_field_type <= _field_stack_stack_num_field_type_16_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h8 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_8_field_type_16_sub_class_id <= _field_stack_stack_num_field_type_16_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h8 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_8_field_type_17_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_17_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h8 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_8_field_type_17_field_type <= _field_stack_stack_num_field_type_17_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h8 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_8_field_type_17_sub_class_id <= _field_stack_stack_num_field_type_17_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h8 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_8_field_type_18_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_18_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h8 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_8_field_type_18_field_type <= _field_stack_stack_num_field_type_18_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h8 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_8_field_type_18_sub_class_id <= _field_stack_stack_num_field_type_18_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h8 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_8_field_type_19_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_19_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h8 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_8_field_type_19_field_type <= _field_stack_stack_num_field_type_19_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h8 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_8_field_type_19_sub_class_id <= _field_stack_stack_num_field_type_19_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h8 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_8_field_type_20_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_20_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h8 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_8_field_type_20_field_type <= _field_stack_stack_num_field_type_20_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h8 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_8_field_type_20_sub_class_id <= _field_stack_stack_num_field_type_20_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h8 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_8_field_type_21_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_21_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h8 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_8_field_type_21_field_type <= _field_stack_stack_num_field_type_21_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h8 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_8_field_type_21_sub_class_id <= _field_stack_stack_num_field_type_21_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h8 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_8_field_type_22_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_22_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h8 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_8_field_type_22_field_type <= _field_stack_stack_num_field_type_22_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h8 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_8_field_type_22_sub_class_id <= _field_stack_stack_num_field_type_22_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h8 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_8_field_type_23_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_23_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h8 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_8_field_type_23_field_type <= _field_stack_stack_num_field_type_23_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h8 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_8_field_type_23_sub_class_id <= _field_stack_stack_num_field_type_23_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h8 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_8_field_type_24_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_24_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h8 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_8_field_type_24_field_type <= _field_stack_stack_num_field_type_24_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h8 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_8_field_type_24_sub_class_id <= _field_stack_stack_num_field_type_24_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h8 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_8_field_type_25_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_25_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h8 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_8_field_type_25_field_type <= _field_stack_stack_num_field_type_25_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h8 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_8_field_type_25_sub_class_id <= _field_stack_stack_num_field_type_25_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h8 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_8_field_type_26_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_26_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h8 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_8_field_type_26_field_type <= _field_stack_stack_num_field_type_26_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h8 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_8_field_type_26_sub_class_id <= _field_stack_stack_num_field_type_26_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h8 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_8_field_type_27_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_27_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h8 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_8_field_type_27_field_type <= _field_stack_stack_num_field_type_27_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h8 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_8_field_type_27_sub_class_id <= _field_stack_stack_num_field_type_27_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h8 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_8_field_type_28_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_28_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h8 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_8_field_type_28_field_type <= _field_stack_stack_num_field_type_28_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h8 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_8_field_type_28_sub_class_id <= _field_stack_stack_num_field_type_28_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h8 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_8_field_type_29_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_29_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h8 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_8_field_type_29_field_type <= _field_stack_stack_num_field_type_29_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h8 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_8_field_type_29_sub_class_id <= _field_stack_stack_num_field_type_29_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h8 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_8_field_type_30_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_30_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h8 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_8_field_type_30_field_type <= _field_stack_stack_num_field_type_30_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h8 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_8_field_type_30_sub_class_id <= _field_stack_stack_num_field_type_30_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h8 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_8_field_type_31_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_31_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h8 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_8_field_type_31_field_type <= _field_stack_stack_num_field_type_31_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h8 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_8_field_type_31_sub_class_id <= _field_stack_stack_num_field_type_31_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h8 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_8_field_type_32_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_32_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h8 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_8_field_type_32_field_type <= _field_stack_stack_num_field_type_32_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h8 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_8_field_type_32_sub_class_id <= _field_stack_stack_num_field_type_32_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h9 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_9_field_type_0_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_0_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h9 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_9_field_type_0_field_type <= _field_stack_stack_num_field_type_0_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h9 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_9_field_type_0_sub_class_id <= _field_stack_stack_num_field_type_0_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h9 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_9_field_type_1_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_1_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h9 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_9_field_type_1_field_type <= _field_stack_stack_num_field_type_1_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h9 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_9_field_type_1_sub_class_id <= _field_stack_stack_num_field_type_1_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h9 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_9_field_type_2_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_2_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h9 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_9_field_type_2_field_type <= _field_stack_stack_num_field_type_2_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h9 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_9_field_type_2_sub_class_id <= _field_stack_stack_num_field_type_2_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h9 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_9_field_type_3_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_3_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h9 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_9_field_type_3_field_type <= _field_stack_stack_num_field_type_3_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h9 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_9_field_type_3_sub_class_id <= _field_stack_stack_num_field_type_3_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h9 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_9_field_type_4_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_4_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h9 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_9_field_type_4_field_type <= _field_stack_stack_num_field_type_4_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h9 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_9_field_type_4_sub_class_id <= _field_stack_stack_num_field_type_4_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h9 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_9_field_type_5_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_5_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h9 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_9_field_type_5_field_type <= _field_stack_stack_num_field_type_5_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h9 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_9_field_type_5_sub_class_id <= _field_stack_stack_num_field_type_5_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h9 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_9_field_type_6_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_6_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h9 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_9_field_type_6_field_type <= _field_stack_stack_num_field_type_6_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h9 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_9_field_type_6_sub_class_id <= _field_stack_stack_num_field_type_6_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h9 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_9_field_type_7_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_7_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h9 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_9_field_type_7_field_type <= _field_stack_stack_num_field_type_7_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h9 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_9_field_type_7_sub_class_id <= _field_stack_stack_num_field_type_7_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h9 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_9_field_type_8_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_8_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h9 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_9_field_type_8_field_type <= _field_stack_stack_num_field_type_8_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h9 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_9_field_type_8_sub_class_id <= _field_stack_stack_num_field_type_8_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h9 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_9_field_type_9_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_9_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h9 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_9_field_type_9_field_type <= _field_stack_stack_num_field_type_9_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h9 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_9_field_type_9_sub_class_id <= _field_stack_stack_num_field_type_9_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h9 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_9_field_type_10_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_10_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h9 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_9_field_type_10_field_type <= _field_stack_stack_num_field_type_10_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h9 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_9_field_type_10_sub_class_id <= _field_stack_stack_num_field_type_10_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h9 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_9_field_type_11_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_11_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h9 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_9_field_type_11_field_type <= _field_stack_stack_num_field_type_11_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h9 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_9_field_type_11_sub_class_id <= _field_stack_stack_num_field_type_11_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h9 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_9_field_type_12_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_12_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h9 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_9_field_type_12_field_type <= _field_stack_stack_num_field_type_12_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h9 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_9_field_type_12_sub_class_id <= _field_stack_stack_num_field_type_12_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h9 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_9_field_type_13_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_13_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h9 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_9_field_type_13_field_type <= _field_stack_stack_num_field_type_13_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h9 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_9_field_type_13_sub_class_id <= _field_stack_stack_num_field_type_13_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h9 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_9_field_type_14_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_14_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h9 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_9_field_type_14_field_type <= _field_stack_stack_num_field_type_14_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h9 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_9_field_type_14_sub_class_id <= _field_stack_stack_num_field_type_14_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h9 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_9_field_type_15_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_15_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h9 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_9_field_type_15_field_type <= _field_stack_stack_num_field_type_15_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h9 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_9_field_type_15_sub_class_id <= _field_stack_stack_num_field_type_15_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h9 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_9_field_type_16_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_16_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h9 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_9_field_type_16_field_type <= _field_stack_stack_num_field_type_16_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h9 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_9_field_type_16_sub_class_id <= _field_stack_stack_num_field_type_16_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h9 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_9_field_type_17_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_17_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h9 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_9_field_type_17_field_type <= _field_stack_stack_num_field_type_17_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h9 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_9_field_type_17_sub_class_id <= _field_stack_stack_num_field_type_17_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h9 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_9_field_type_18_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_18_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h9 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_9_field_type_18_field_type <= _field_stack_stack_num_field_type_18_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h9 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_9_field_type_18_sub_class_id <= _field_stack_stack_num_field_type_18_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h9 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_9_field_type_19_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_19_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h9 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_9_field_type_19_field_type <= _field_stack_stack_num_field_type_19_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h9 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_9_field_type_19_sub_class_id <= _field_stack_stack_num_field_type_19_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h9 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_9_field_type_20_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_20_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h9 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_9_field_type_20_field_type <= _field_stack_stack_num_field_type_20_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h9 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_9_field_type_20_sub_class_id <= _field_stack_stack_num_field_type_20_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h9 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_9_field_type_21_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_21_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h9 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_9_field_type_21_field_type <= _field_stack_stack_num_field_type_21_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h9 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_9_field_type_21_sub_class_id <= _field_stack_stack_num_field_type_21_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h9 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_9_field_type_22_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_22_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h9 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_9_field_type_22_field_type <= _field_stack_stack_num_field_type_22_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h9 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_9_field_type_22_sub_class_id <= _field_stack_stack_num_field_type_22_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h9 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_9_field_type_23_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_23_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h9 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_9_field_type_23_field_type <= _field_stack_stack_num_field_type_23_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h9 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_9_field_type_23_sub_class_id <= _field_stack_stack_num_field_type_23_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h9 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_9_field_type_24_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_24_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h9 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_9_field_type_24_field_type <= _field_stack_stack_num_field_type_24_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h9 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_9_field_type_24_sub_class_id <= _field_stack_stack_num_field_type_24_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h9 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_9_field_type_25_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_25_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h9 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_9_field_type_25_field_type <= _field_stack_stack_num_field_type_25_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h9 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_9_field_type_25_sub_class_id <= _field_stack_stack_num_field_type_25_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h9 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_9_field_type_26_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_26_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h9 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_9_field_type_26_field_type <= _field_stack_stack_num_field_type_26_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h9 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_9_field_type_26_sub_class_id <= _field_stack_stack_num_field_type_26_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h9 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_9_field_type_27_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_27_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h9 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_9_field_type_27_field_type <= _field_stack_stack_num_field_type_27_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h9 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_9_field_type_27_sub_class_id <= _field_stack_stack_num_field_type_27_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h9 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_9_field_type_28_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_28_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h9 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_9_field_type_28_field_type <= _field_stack_stack_num_field_type_28_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h9 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_9_field_type_28_sub_class_id <= _field_stack_stack_num_field_type_28_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h9 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_9_field_type_29_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_29_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h9 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_9_field_type_29_field_type <= _field_stack_stack_num_field_type_29_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h9 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_9_field_type_29_sub_class_id <= _field_stack_stack_num_field_type_29_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h9 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_9_field_type_30_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_30_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h9 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_9_field_type_30_field_type <= _field_stack_stack_num_field_type_30_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h9 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_9_field_type_30_sub_class_id <= _field_stack_stack_num_field_type_30_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h9 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_9_field_type_31_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_31_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h9 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_9_field_type_31_field_type <= _field_stack_stack_num_field_type_31_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h9 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_9_field_type_31_sub_class_id <= _field_stack_stack_num_field_type_31_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h9 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_9_field_type_32_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_32_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h9 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_9_field_type_32_field_type <= _field_stack_stack_num_field_type_32_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'h9 == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_9_field_type_32_sub_class_id <= _field_stack_stack_num_field_type_32_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'ha == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_10_field_type_0_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_0_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'ha == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_10_field_type_0_field_type <= _field_stack_stack_num_field_type_0_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'ha == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_10_field_type_0_sub_class_id <= _field_stack_stack_num_field_type_0_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'ha == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_10_field_type_1_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_1_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'ha == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_10_field_type_1_field_type <= _field_stack_stack_num_field_type_1_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'ha == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_10_field_type_1_sub_class_id <= _field_stack_stack_num_field_type_1_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'ha == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_10_field_type_2_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_2_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'ha == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_10_field_type_2_field_type <= _field_stack_stack_num_field_type_2_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'ha == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_10_field_type_2_sub_class_id <= _field_stack_stack_num_field_type_2_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'ha == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_10_field_type_3_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_3_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'ha == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_10_field_type_3_field_type <= _field_stack_stack_num_field_type_3_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'ha == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_10_field_type_3_sub_class_id <= _field_stack_stack_num_field_type_3_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'ha == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_10_field_type_4_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_4_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'ha == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_10_field_type_4_field_type <= _field_stack_stack_num_field_type_4_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'ha == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_10_field_type_4_sub_class_id <= _field_stack_stack_num_field_type_4_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'ha == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_10_field_type_5_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_5_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'ha == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_10_field_type_5_field_type <= _field_stack_stack_num_field_type_5_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'ha == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_10_field_type_5_sub_class_id <= _field_stack_stack_num_field_type_5_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'ha == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_10_field_type_6_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_6_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'ha == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_10_field_type_6_field_type <= _field_stack_stack_num_field_type_6_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'ha == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_10_field_type_6_sub_class_id <= _field_stack_stack_num_field_type_6_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'ha == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_10_field_type_7_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_7_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'ha == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_10_field_type_7_field_type <= _field_stack_stack_num_field_type_7_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'ha == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_10_field_type_7_sub_class_id <= _field_stack_stack_num_field_type_7_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'ha == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_10_field_type_8_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_8_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'ha == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_10_field_type_8_field_type <= _field_stack_stack_num_field_type_8_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'ha == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_10_field_type_8_sub_class_id <= _field_stack_stack_num_field_type_8_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'ha == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_10_field_type_9_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_9_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'ha == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_10_field_type_9_field_type <= _field_stack_stack_num_field_type_9_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'ha == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_10_field_type_9_sub_class_id <= _field_stack_stack_num_field_type_9_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'ha == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_10_field_type_10_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_10_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'ha == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_10_field_type_10_field_type <= _field_stack_stack_num_field_type_10_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'ha == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_10_field_type_10_sub_class_id <= _field_stack_stack_num_field_type_10_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'ha == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_10_field_type_11_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_11_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'ha == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_10_field_type_11_field_type <= _field_stack_stack_num_field_type_11_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'ha == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_10_field_type_11_sub_class_id <= _field_stack_stack_num_field_type_11_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'ha == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_10_field_type_12_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_12_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'ha == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_10_field_type_12_field_type <= _field_stack_stack_num_field_type_12_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'ha == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_10_field_type_12_sub_class_id <= _field_stack_stack_num_field_type_12_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'ha == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_10_field_type_13_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_13_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'ha == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_10_field_type_13_field_type <= _field_stack_stack_num_field_type_13_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'ha == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_10_field_type_13_sub_class_id <= _field_stack_stack_num_field_type_13_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'ha == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_10_field_type_14_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_14_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'ha == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_10_field_type_14_field_type <= _field_stack_stack_num_field_type_14_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'ha == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_10_field_type_14_sub_class_id <= _field_stack_stack_num_field_type_14_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'ha == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_10_field_type_15_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_15_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'ha == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_10_field_type_15_field_type <= _field_stack_stack_num_field_type_15_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'ha == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_10_field_type_15_sub_class_id <= _field_stack_stack_num_field_type_15_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'ha == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_10_field_type_16_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_16_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'ha == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_10_field_type_16_field_type <= _field_stack_stack_num_field_type_16_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'ha == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_10_field_type_16_sub_class_id <= _field_stack_stack_num_field_type_16_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'ha == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_10_field_type_17_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_17_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'ha == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_10_field_type_17_field_type <= _field_stack_stack_num_field_type_17_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'ha == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_10_field_type_17_sub_class_id <= _field_stack_stack_num_field_type_17_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'ha == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_10_field_type_18_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_18_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'ha == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_10_field_type_18_field_type <= _field_stack_stack_num_field_type_18_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'ha == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_10_field_type_18_sub_class_id <= _field_stack_stack_num_field_type_18_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'ha == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_10_field_type_19_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_19_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'ha == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_10_field_type_19_field_type <= _field_stack_stack_num_field_type_19_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'ha == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_10_field_type_19_sub_class_id <= _field_stack_stack_num_field_type_19_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'ha == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_10_field_type_20_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_20_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'ha == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_10_field_type_20_field_type <= _field_stack_stack_num_field_type_20_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'ha == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_10_field_type_20_sub_class_id <= _field_stack_stack_num_field_type_20_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'ha == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_10_field_type_21_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_21_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'ha == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_10_field_type_21_field_type <= _field_stack_stack_num_field_type_21_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'ha == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_10_field_type_21_sub_class_id <= _field_stack_stack_num_field_type_21_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'ha == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_10_field_type_22_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_22_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'ha == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_10_field_type_22_field_type <= _field_stack_stack_num_field_type_22_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'ha == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_10_field_type_22_sub_class_id <= _field_stack_stack_num_field_type_22_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'ha == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_10_field_type_23_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_23_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'ha == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_10_field_type_23_field_type <= _field_stack_stack_num_field_type_23_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'ha == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_10_field_type_23_sub_class_id <= _field_stack_stack_num_field_type_23_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'ha == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_10_field_type_24_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_24_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'ha == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_10_field_type_24_field_type <= _field_stack_stack_num_field_type_24_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'ha == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_10_field_type_24_sub_class_id <= _field_stack_stack_num_field_type_24_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'ha == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_10_field_type_25_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_25_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'ha == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_10_field_type_25_field_type <= _field_stack_stack_num_field_type_25_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'ha == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_10_field_type_25_sub_class_id <= _field_stack_stack_num_field_type_25_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'ha == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_10_field_type_26_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_26_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'ha == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_10_field_type_26_field_type <= _field_stack_stack_num_field_type_26_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'ha == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_10_field_type_26_sub_class_id <= _field_stack_stack_num_field_type_26_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'ha == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_10_field_type_27_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_27_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'ha == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_10_field_type_27_field_type <= _field_stack_stack_num_field_type_27_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'ha == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_10_field_type_27_sub_class_id <= _field_stack_stack_num_field_type_27_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'ha == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_10_field_type_28_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_28_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'ha == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_10_field_type_28_field_type <= _field_stack_stack_num_field_type_28_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'ha == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_10_field_type_28_sub_class_id <= _field_stack_stack_num_field_type_28_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'ha == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_10_field_type_29_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_29_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'ha == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_10_field_type_29_field_type <= _field_stack_stack_num_field_type_29_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'ha == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_10_field_type_29_sub_class_id <= _field_stack_stack_num_field_type_29_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'ha == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_10_field_type_30_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_30_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'ha == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_10_field_type_30_field_type <= _field_stack_stack_num_field_type_30_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'ha == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_10_field_type_30_sub_class_id <= _field_stack_stack_num_field_type_30_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'ha == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_10_field_type_31_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_31_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'ha == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_10_field_type_31_field_type <= _field_stack_stack_num_field_type_31_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'ha == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_10_field_type_31_sub_class_id <= _field_stack_stack_num_field_type_31_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'ha == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_10_field_type_32_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_32_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'ha == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_10_field_type_32_field_type <= _field_stack_stack_num_field_type_32_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'ha == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_10_field_type_32_sub_class_id <= _field_stack_stack_num_field_type_32_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hb == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_11_field_type_0_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_0_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hb == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_11_field_type_0_field_type <= _field_stack_stack_num_field_type_0_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hb == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_11_field_type_0_sub_class_id <= _field_stack_stack_num_field_type_0_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hb == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_11_field_type_1_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_1_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hb == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_11_field_type_1_field_type <= _field_stack_stack_num_field_type_1_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hb == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_11_field_type_1_sub_class_id <= _field_stack_stack_num_field_type_1_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hb == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_11_field_type_2_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_2_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hb == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_11_field_type_2_field_type <= _field_stack_stack_num_field_type_2_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hb == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_11_field_type_2_sub_class_id <= _field_stack_stack_num_field_type_2_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hb == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_11_field_type_3_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_3_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hb == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_11_field_type_3_field_type <= _field_stack_stack_num_field_type_3_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hb == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_11_field_type_3_sub_class_id <= _field_stack_stack_num_field_type_3_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hb == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_11_field_type_4_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_4_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hb == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_11_field_type_4_field_type <= _field_stack_stack_num_field_type_4_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hb == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_11_field_type_4_sub_class_id <= _field_stack_stack_num_field_type_4_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hb == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_11_field_type_5_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_5_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hb == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_11_field_type_5_field_type <= _field_stack_stack_num_field_type_5_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hb == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_11_field_type_5_sub_class_id <= _field_stack_stack_num_field_type_5_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hb == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_11_field_type_6_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_6_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hb == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_11_field_type_6_field_type <= _field_stack_stack_num_field_type_6_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hb == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_11_field_type_6_sub_class_id <= _field_stack_stack_num_field_type_6_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hb == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_11_field_type_7_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_7_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hb == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_11_field_type_7_field_type <= _field_stack_stack_num_field_type_7_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hb == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_11_field_type_7_sub_class_id <= _field_stack_stack_num_field_type_7_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hb == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_11_field_type_8_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_8_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hb == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_11_field_type_8_field_type <= _field_stack_stack_num_field_type_8_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hb == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_11_field_type_8_sub_class_id <= _field_stack_stack_num_field_type_8_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hb == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_11_field_type_9_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_9_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hb == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_11_field_type_9_field_type <= _field_stack_stack_num_field_type_9_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hb == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_11_field_type_9_sub_class_id <= _field_stack_stack_num_field_type_9_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hb == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_11_field_type_10_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_10_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hb == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_11_field_type_10_field_type <= _field_stack_stack_num_field_type_10_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hb == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_11_field_type_10_sub_class_id <= _field_stack_stack_num_field_type_10_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hb == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_11_field_type_11_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_11_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hb == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_11_field_type_11_field_type <= _field_stack_stack_num_field_type_11_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hb == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_11_field_type_11_sub_class_id <= _field_stack_stack_num_field_type_11_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hb == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_11_field_type_12_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_12_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hb == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_11_field_type_12_field_type <= _field_stack_stack_num_field_type_12_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hb == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_11_field_type_12_sub_class_id <= _field_stack_stack_num_field_type_12_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hb == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_11_field_type_13_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_13_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hb == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_11_field_type_13_field_type <= _field_stack_stack_num_field_type_13_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hb == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_11_field_type_13_sub_class_id <= _field_stack_stack_num_field_type_13_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hb == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_11_field_type_14_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_14_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hb == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_11_field_type_14_field_type <= _field_stack_stack_num_field_type_14_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hb == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_11_field_type_14_sub_class_id <= _field_stack_stack_num_field_type_14_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hb == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_11_field_type_15_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_15_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hb == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_11_field_type_15_field_type <= _field_stack_stack_num_field_type_15_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hb == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_11_field_type_15_sub_class_id <= _field_stack_stack_num_field_type_15_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hb == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_11_field_type_16_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_16_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hb == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_11_field_type_16_field_type <= _field_stack_stack_num_field_type_16_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hb == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_11_field_type_16_sub_class_id <= _field_stack_stack_num_field_type_16_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hb == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_11_field_type_17_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_17_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hb == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_11_field_type_17_field_type <= _field_stack_stack_num_field_type_17_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hb == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_11_field_type_17_sub_class_id <= _field_stack_stack_num_field_type_17_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hb == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_11_field_type_18_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_18_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hb == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_11_field_type_18_field_type <= _field_stack_stack_num_field_type_18_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hb == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_11_field_type_18_sub_class_id <= _field_stack_stack_num_field_type_18_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hb == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_11_field_type_19_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_19_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hb == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_11_field_type_19_field_type <= _field_stack_stack_num_field_type_19_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hb == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_11_field_type_19_sub_class_id <= _field_stack_stack_num_field_type_19_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hb == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_11_field_type_20_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_20_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hb == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_11_field_type_20_field_type <= _field_stack_stack_num_field_type_20_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hb == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_11_field_type_20_sub_class_id <= _field_stack_stack_num_field_type_20_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hb == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_11_field_type_21_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_21_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hb == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_11_field_type_21_field_type <= _field_stack_stack_num_field_type_21_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hb == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_11_field_type_21_sub_class_id <= _field_stack_stack_num_field_type_21_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hb == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_11_field_type_22_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_22_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hb == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_11_field_type_22_field_type <= _field_stack_stack_num_field_type_22_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hb == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_11_field_type_22_sub_class_id <= _field_stack_stack_num_field_type_22_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hb == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_11_field_type_23_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_23_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hb == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_11_field_type_23_field_type <= _field_stack_stack_num_field_type_23_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hb == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_11_field_type_23_sub_class_id <= _field_stack_stack_num_field_type_23_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hb == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_11_field_type_24_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_24_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hb == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_11_field_type_24_field_type <= _field_stack_stack_num_field_type_24_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hb == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_11_field_type_24_sub_class_id <= _field_stack_stack_num_field_type_24_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hb == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_11_field_type_25_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_25_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hb == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_11_field_type_25_field_type <= _field_stack_stack_num_field_type_25_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hb == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_11_field_type_25_sub_class_id <= _field_stack_stack_num_field_type_25_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hb == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_11_field_type_26_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_26_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hb == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_11_field_type_26_field_type <= _field_stack_stack_num_field_type_26_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hb == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_11_field_type_26_sub_class_id <= _field_stack_stack_num_field_type_26_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hb == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_11_field_type_27_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_27_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hb == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_11_field_type_27_field_type <= _field_stack_stack_num_field_type_27_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hb == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_11_field_type_27_sub_class_id <= _field_stack_stack_num_field_type_27_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hb == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_11_field_type_28_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_28_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hb == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_11_field_type_28_field_type <= _field_stack_stack_num_field_type_28_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hb == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_11_field_type_28_sub_class_id <= _field_stack_stack_num_field_type_28_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hb == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_11_field_type_29_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_29_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hb == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_11_field_type_29_field_type <= _field_stack_stack_num_field_type_29_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hb == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_11_field_type_29_sub_class_id <= _field_stack_stack_num_field_type_29_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hb == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_11_field_type_30_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_30_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hb == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_11_field_type_30_field_type <= _field_stack_stack_num_field_type_30_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hb == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_11_field_type_30_sub_class_id <= _field_stack_stack_num_field_type_30_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hb == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_11_field_type_31_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_31_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hb == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_11_field_type_31_field_type <= _field_stack_stack_num_field_type_31_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hb == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_11_field_type_31_sub_class_id <= _field_stack_stack_num_field_type_31_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hb == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_11_field_type_32_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_32_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hb == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_11_field_type_32_field_type <= _field_stack_stack_num_field_type_32_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hb == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_11_field_type_32_sub_class_id <= _field_stack_stack_num_field_type_32_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hc == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_12_field_type_0_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_0_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hc == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_12_field_type_0_field_type <= _field_stack_stack_num_field_type_0_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hc == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_12_field_type_0_sub_class_id <= _field_stack_stack_num_field_type_0_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hc == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_12_field_type_1_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_1_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hc == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_12_field_type_1_field_type <= _field_stack_stack_num_field_type_1_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hc == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_12_field_type_1_sub_class_id <= _field_stack_stack_num_field_type_1_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hc == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_12_field_type_2_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_2_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hc == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_12_field_type_2_field_type <= _field_stack_stack_num_field_type_2_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hc == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_12_field_type_2_sub_class_id <= _field_stack_stack_num_field_type_2_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hc == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_12_field_type_3_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_3_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hc == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_12_field_type_3_field_type <= _field_stack_stack_num_field_type_3_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hc == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_12_field_type_3_sub_class_id <= _field_stack_stack_num_field_type_3_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hc == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_12_field_type_4_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_4_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hc == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_12_field_type_4_field_type <= _field_stack_stack_num_field_type_4_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hc == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_12_field_type_4_sub_class_id <= _field_stack_stack_num_field_type_4_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hc == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_12_field_type_5_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_5_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hc == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_12_field_type_5_field_type <= _field_stack_stack_num_field_type_5_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hc == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_12_field_type_5_sub_class_id <= _field_stack_stack_num_field_type_5_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hc == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_12_field_type_6_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_6_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hc == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_12_field_type_6_field_type <= _field_stack_stack_num_field_type_6_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hc == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_12_field_type_6_sub_class_id <= _field_stack_stack_num_field_type_6_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hc == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_12_field_type_7_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_7_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hc == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_12_field_type_7_field_type <= _field_stack_stack_num_field_type_7_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hc == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_12_field_type_7_sub_class_id <= _field_stack_stack_num_field_type_7_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hc == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_12_field_type_8_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_8_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hc == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_12_field_type_8_field_type <= _field_stack_stack_num_field_type_8_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hc == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_12_field_type_8_sub_class_id <= _field_stack_stack_num_field_type_8_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hc == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_12_field_type_9_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_9_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hc == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_12_field_type_9_field_type <= _field_stack_stack_num_field_type_9_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hc == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_12_field_type_9_sub_class_id <= _field_stack_stack_num_field_type_9_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hc == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_12_field_type_10_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_10_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hc == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_12_field_type_10_field_type <= _field_stack_stack_num_field_type_10_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hc == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_12_field_type_10_sub_class_id <= _field_stack_stack_num_field_type_10_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hc == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_12_field_type_11_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_11_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hc == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_12_field_type_11_field_type <= _field_stack_stack_num_field_type_11_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hc == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_12_field_type_11_sub_class_id <= _field_stack_stack_num_field_type_11_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hc == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_12_field_type_12_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_12_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hc == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_12_field_type_12_field_type <= _field_stack_stack_num_field_type_12_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hc == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_12_field_type_12_sub_class_id <= _field_stack_stack_num_field_type_12_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hc == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_12_field_type_13_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_13_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hc == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_12_field_type_13_field_type <= _field_stack_stack_num_field_type_13_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hc == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_12_field_type_13_sub_class_id <= _field_stack_stack_num_field_type_13_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hc == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_12_field_type_14_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_14_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hc == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_12_field_type_14_field_type <= _field_stack_stack_num_field_type_14_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hc == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_12_field_type_14_sub_class_id <= _field_stack_stack_num_field_type_14_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hc == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_12_field_type_15_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_15_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hc == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_12_field_type_15_field_type <= _field_stack_stack_num_field_type_15_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hc == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_12_field_type_15_sub_class_id <= _field_stack_stack_num_field_type_15_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hc == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_12_field_type_16_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_16_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hc == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_12_field_type_16_field_type <= _field_stack_stack_num_field_type_16_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hc == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_12_field_type_16_sub_class_id <= _field_stack_stack_num_field_type_16_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hc == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_12_field_type_17_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_17_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hc == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_12_field_type_17_field_type <= _field_stack_stack_num_field_type_17_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hc == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_12_field_type_17_sub_class_id <= _field_stack_stack_num_field_type_17_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hc == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_12_field_type_18_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_18_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hc == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_12_field_type_18_field_type <= _field_stack_stack_num_field_type_18_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hc == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_12_field_type_18_sub_class_id <= _field_stack_stack_num_field_type_18_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hc == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_12_field_type_19_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_19_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hc == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_12_field_type_19_field_type <= _field_stack_stack_num_field_type_19_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hc == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_12_field_type_19_sub_class_id <= _field_stack_stack_num_field_type_19_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hc == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_12_field_type_20_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_20_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hc == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_12_field_type_20_field_type <= _field_stack_stack_num_field_type_20_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hc == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_12_field_type_20_sub_class_id <= _field_stack_stack_num_field_type_20_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hc == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_12_field_type_21_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_21_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hc == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_12_field_type_21_field_type <= _field_stack_stack_num_field_type_21_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hc == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_12_field_type_21_sub_class_id <= _field_stack_stack_num_field_type_21_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hc == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_12_field_type_22_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_22_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hc == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_12_field_type_22_field_type <= _field_stack_stack_num_field_type_22_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hc == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_12_field_type_22_sub_class_id <= _field_stack_stack_num_field_type_22_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hc == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_12_field_type_23_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_23_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hc == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_12_field_type_23_field_type <= _field_stack_stack_num_field_type_23_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hc == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_12_field_type_23_sub_class_id <= _field_stack_stack_num_field_type_23_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hc == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_12_field_type_24_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_24_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hc == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_12_field_type_24_field_type <= _field_stack_stack_num_field_type_24_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hc == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_12_field_type_24_sub_class_id <= _field_stack_stack_num_field_type_24_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hc == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_12_field_type_25_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_25_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hc == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_12_field_type_25_field_type <= _field_stack_stack_num_field_type_25_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hc == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_12_field_type_25_sub_class_id <= _field_stack_stack_num_field_type_25_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hc == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_12_field_type_26_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_26_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hc == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_12_field_type_26_field_type <= _field_stack_stack_num_field_type_26_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hc == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_12_field_type_26_sub_class_id <= _field_stack_stack_num_field_type_26_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hc == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_12_field_type_27_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_27_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hc == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_12_field_type_27_field_type <= _field_stack_stack_num_field_type_27_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hc == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_12_field_type_27_sub_class_id <= _field_stack_stack_num_field_type_27_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hc == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_12_field_type_28_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_28_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hc == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_12_field_type_28_field_type <= _field_stack_stack_num_field_type_28_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hc == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_12_field_type_28_sub_class_id <= _field_stack_stack_num_field_type_28_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hc == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_12_field_type_29_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_29_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hc == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_12_field_type_29_field_type <= _field_stack_stack_num_field_type_29_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hc == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_12_field_type_29_sub_class_id <= _field_stack_stack_num_field_type_29_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hc == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_12_field_type_30_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_30_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hc == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_12_field_type_30_field_type <= _field_stack_stack_num_field_type_30_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hc == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_12_field_type_30_sub_class_id <= _field_stack_stack_num_field_type_30_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hc == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_12_field_type_31_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_31_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hc == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_12_field_type_31_field_type <= _field_stack_stack_num_field_type_31_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hc == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_12_field_type_31_sub_class_id <= _field_stack_stack_num_field_type_31_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hc == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_12_field_type_32_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_32_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hc == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_12_field_type_32_field_type <= _field_stack_stack_num_field_type_32_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hc == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_12_field_type_32_sub_class_id <= _field_stack_stack_num_field_type_32_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hd == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_13_field_type_0_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_0_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hd == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_13_field_type_0_field_type <= _field_stack_stack_num_field_type_0_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hd == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_13_field_type_0_sub_class_id <= _field_stack_stack_num_field_type_0_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hd == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_13_field_type_1_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_1_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hd == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_13_field_type_1_field_type <= _field_stack_stack_num_field_type_1_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hd == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_13_field_type_1_sub_class_id <= _field_stack_stack_num_field_type_1_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hd == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_13_field_type_2_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_2_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hd == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_13_field_type_2_field_type <= _field_stack_stack_num_field_type_2_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hd == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_13_field_type_2_sub_class_id <= _field_stack_stack_num_field_type_2_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hd == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_13_field_type_3_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_3_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hd == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_13_field_type_3_field_type <= _field_stack_stack_num_field_type_3_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hd == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_13_field_type_3_sub_class_id <= _field_stack_stack_num_field_type_3_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hd == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_13_field_type_4_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_4_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hd == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_13_field_type_4_field_type <= _field_stack_stack_num_field_type_4_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hd == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_13_field_type_4_sub_class_id <= _field_stack_stack_num_field_type_4_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hd == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_13_field_type_5_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_5_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hd == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_13_field_type_5_field_type <= _field_stack_stack_num_field_type_5_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hd == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_13_field_type_5_sub_class_id <= _field_stack_stack_num_field_type_5_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hd == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_13_field_type_6_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_6_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hd == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_13_field_type_6_field_type <= _field_stack_stack_num_field_type_6_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hd == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_13_field_type_6_sub_class_id <= _field_stack_stack_num_field_type_6_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hd == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_13_field_type_7_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_7_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hd == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_13_field_type_7_field_type <= _field_stack_stack_num_field_type_7_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hd == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_13_field_type_7_sub_class_id <= _field_stack_stack_num_field_type_7_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hd == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_13_field_type_8_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_8_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hd == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_13_field_type_8_field_type <= _field_stack_stack_num_field_type_8_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hd == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_13_field_type_8_sub_class_id <= _field_stack_stack_num_field_type_8_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hd == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_13_field_type_9_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_9_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hd == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_13_field_type_9_field_type <= _field_stack_stack_num_field_type_9_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hd == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_13_field_type_9_sub_class_id <= _field_stack_stack_num_field_type_9_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hd == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_13_field_type_10_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_10_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hd == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_13_field_type_10_field_type <= _field_stack_stack_num_field_type_10_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hd == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_13_field_type_10_sub_class_id <= _field_stack_stack_num_field_type_10_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hd == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_13_field_type_11_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_11_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hd == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_13_field_type_11_field_type <= _field_stack_stack_num_field_type_11_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hd == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_13_field_type_11_sub_class_id <= _field_stack_stack_num_field_type_11_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hd == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_13_field_type_12_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_12_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hd == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_13_field_type_12_field_type <= _field_stack_stack_num_field_type_12_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hd == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_13_field_type_12_sub_class_id <= _field_stack_stack_num_field_type_12_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hd == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_13_field_type_13_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_13_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hd == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_13_field_type_13_field_type <= _field_stack_stack_num_field_type_13_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hd == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_13_field_type_13_sub_class_id <= _field_stack_stack_num_field_type_13_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hd == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_13_field_type_14_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_14_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hd == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_13_field_type_14_field_type <= _field_stack_stack_num_field_type_14_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hd == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_13_field_type_14_sub_class_id <= _field_stack_stack_num_field_type_14_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hd == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_13_field_type_15_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_15_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hd == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_13_field_type_15_field_type <= _field_stack_stack_num_field_type_15_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hd == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_13_field_type_15_sub_class_id <= _field_stack_stack_num_field_type_15_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hd == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_13_field_type_16_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_16_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hd == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_13_field_type_16_field_type <= _field_stack_stack_num_field_type_16_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hd == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_13_field_type_16_sub_class_id <= _field_stack_stack_num_field_type_16_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hd == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_13_field_type_17_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_17_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hd == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_13_field_type_17_field_type <= _field_stack_stack_num_field_type_17_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hd == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_13_field_type_17_sub_class_id <= _field_stack_stack_num_field_type_17_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hd == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_13_field_type_18_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_18_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hd == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_13_field_type_18_field_type <= _field_stack_stack_num_field_type_18_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hd == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_13_field_type_18_sub_class_id <= _field_stack_stack_num_field_type_18_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hd == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_13_field_type_19_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_19_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hd == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_13_field_type_19_field_type <= _field_stack_stack_num_field_type_19_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hd == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_13_field_type_19_sub_class_id <= _field_stack_stack_num_field_type_19_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hd == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_13_field_type_20_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_20_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hd == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_13_field_type_20_field_type <= _field_stack_stack_num_field_type_20_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hd == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_13_field_type_20_sub_class_id <= _field_stack_stack_num_field_type_20_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hd == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_13_field_type_21_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_21_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hd == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_13_field_type_21_field_type <= _field_stack_stack_num_field_type_21_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hd == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_13_field_type_21_sub_class_id <= _field_stack_stack_num_field_type_21_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hd == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_13_field_type_22_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_22_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hd == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_13_field_type_22_field_type <= _field_stack_stack_num_field_type_22_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hd == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_13_field_type_22_sub_class_id <= _field_stack_stack_num_field_type_22_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hd == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_13_field_type_23_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_23_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hd == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_13_field_type_23_field_type <= _field_stack_stack_num_field_type_23_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hd == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_13_field_type_23_sub_class_id <= _field_stack_stack_num_field_type_23_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hd == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_13_field_type_24_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_24_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hd == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_13_field_type_24_field_type <= _field_stack_stack_num_field_type_24_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hd == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_13_field_type_24_sub_class_id <= _field_stack_stack_num_field_type_24_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hd == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_13_field_type_25_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_25_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hd == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_13_field_type_25_field_type <= _field_stack_stack_num_field_type_25_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hd == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_13_field_type_25_sub_class_id <= _field_stack_stack_num_field_type_25_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hd == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_13_field_type_26_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_26_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hd == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_13_field_type_26_field_type <= _field_stack_stack_num_field_type_26_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hd == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_13_field_type_26_sub_class_id <= _field_stack_stack_num_field_type_26_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hd == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_13_field_type_27_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_27_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hd == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_13_field_type_27_field_type <= _field_stack_stack_num_field_type_27_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hd == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_13_field_type_27_sub_class_id <= _field_stack_stack_num_field_type_27_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hd == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_13_field_type_28_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_28_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hd == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_13_field_type_28_field_type <= _field_stack_stack_num_field_type_28_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hd == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_13_field_type_28_sub_class_id <= _field_stack_stack_num_field_type_28_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hd == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_13_field_type_29_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_29_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hd == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_13_field_type_29_field_type <= _field_stack_stack_num_field_type_29_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hd == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_13_field_type_29_sub_class_id <= _field_stack_stack_num_field_type_29_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hd == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_13_field_type_30_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_30_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hd == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_13_field_type_30_field_type <= _field_stack_stack_num_field_type_30_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hd == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_13_field_type_30_sub_class_id <= _field_stack_stack_num_field_type_30_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hd == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_13_field_type_31_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_31_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hd == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_13_field_type_31_field_type <= _field_stack_stack_num_field_type_31_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hd == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_13_field_type_31_sub_class_id <= _field_stack_stack_num_field_type_31_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hd == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_13_field_type_32_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_32_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hd == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_13_field_type_32_field_type <= _field_stack_stack_num_field_type_32_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'hd == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_13_field_type_32_sub_class_id <= _field_stack_stack_num_field_type_32_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'he == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_14_field_type_0_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_0_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'he == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_14_field_type_0_field_type <= _field_stack_stack_num_field_type_0_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'he == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_14_field_type_0_sub_class_id <= _field_stack_stack_num_field_type_0_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'he == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_14_field_type_1_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_1_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'he == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_14_field_type_1_field_type <= _field_stack_stack_num_field_type_1_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'he == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_14_field_type_1_sub_class_id <= _field_stack_stack_num_field_type_1_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'he == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_14_field_type_2_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_2_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'he == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_14_field_type_2_field_type <= _field_stack_stack_num_field_type_2_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'he == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_14_field_type_2_sub_class_id <= _field_stack_stack_num_field_type_2_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'he == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_14_field_type_3_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_3_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'he == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_14_field_type_3_field_type <= _field_stack_stack_num_field_type_3_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'he == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_14_field_type_3_sub_class_id <= _field_stack_stack_num_field_type_3_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'he == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_14_field_type_4_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_4_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'he == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_14_field_type_4_field_type <= _field_stack_stack_num_field_type_4_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'he == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_14_field_type_4_sub_class_id <= _field_stack_stack_num_field_type_4_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'he == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_14_field_type_5_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_5_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'he == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_14_field_type_5_field_type <= _field_stack_stack_num_field_type_5_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'he == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_14_field_type_5_sub_class_id <= _field_stack_stack_num_field_type_5_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'he == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_14_field_type_6_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_6_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'he == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_14_field_type_6_field_type <= _field_stack_stack_num_field_type_6_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'he == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_14_field_type_6_sub_class_id <= _field_stack_stack_num_field_type_6_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'he == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_14_field_type_7_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_7_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'he == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_14_field_type_7_field_type <= _field_stack_stack_num_field_type_7_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'he == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_14_field_type_7_sub_class_id <= _field_stack_stack_num_field_type_7_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'he == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_14_field_type_8_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_8_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'he == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_14_field_type_8_field_type <= _field_stack_stack_num_field_type_8_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'he == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_14_field_type_8_sub_class_id <= _field_stack_stack_num_field_type_8_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'he == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_14_field_type_9_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_9_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'he == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_14_field_type_9_field_type <= _field_stack_stack_num_field_type_9_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'he == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_14_field_type_9_sub_class_id <= _field_stack_stack_num_field_type_9_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'he == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_14_field_type_10_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_10_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'he == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_14_field_type_10_field_type <= _field_stack_stack_num_field_type_10_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'he == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_14_field_type_10_sub_class_id <= _field_stack_stack_num_field_type_10_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'he == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_14_field_type_11_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_11_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'he == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_14_field_type_11_field_type <= _field_stack_stack_num_field_type_11_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'he == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_14_field_type_11_sub_class_id <= _field_stack_stack_num_field_type_11_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'he == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_14_field_type_12_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_12_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'he == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_14_field_type_12_field_type <= _field_stack_stack_num_field_type_12_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'he == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_14_field_type_12_sub_class_id <= _field_stack_stack_num_field_type_12_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'he == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_14_field_type_13_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_13_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'he == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_14_field_type_13_field_type <= _field_stack_stack_num_field_type_13_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'he == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_14_field_type_13_sub_class_id <= _field_stack_stack_num_field_type_13_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'he == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_14_field_type_14_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_14_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'he == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_14_field_type_14_field_type <= _field_stack_stack_num_field_type_14_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'he == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_14_field_type_14_sub_class_id <= _field_stack_stack_num_field_type_14_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'he == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_14_field_type_15_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_15_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'he == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_14_field_type_15_field_type <= _field_stack_stack_num_field_type_15_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'he == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_14_field_type_15_sub_class_id <= _field_stack_stack_num_field_type_15_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'he == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_14_field_type_16_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_16_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'he == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_14_field_type_16_field_type <= _field_stack_stack_num_field_type_16_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'he == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_14_field_type_16_sub_class_id <= _field_stack_stack_num_field_type_16_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'he == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_14_field_type_17_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_17_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'he == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_14_field_type_17_field_type <= _field_stack_stack_num_field_type_17_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'he == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_14_field_type_17_sub_class_id <= _field_stack_stack_num_field_type_17_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'he == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_14_field_type_18_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_18_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'he == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_14_field_type_18_field_type <= _field_stack_stack_num_field_type_18_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'he == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_14_field_type_18_sub_class_id <= _field_stack_stack_num_field_type_18_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'he == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_14_field_type_19_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_19_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'he == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_14_field_type_19_field_type <= _field_stack_stack_num_field_type_19_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'he == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_14_field_type_19_sub_class_id <= _field_stack_stack_num_field_type_19_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'he == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_14_field_type_20_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_20_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'he == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_14_field_type_20_field_type <= _field_stack_stack_num_field_type_20_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'he == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_14_field_type_20_sub_class_id <= _field_stack_stack_num_field_type_20_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'he == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_14_field_type_21_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_21_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'he == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_14_field_type_21_field_type <= _field_stack_stack_num_field_type_21_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'he == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_14_field_type_21_sub_class_id <= _field_stack_stack_num_field_type_21_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'he == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_14_field_type_22_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_22_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'he == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_14_field_type_22_field_type <= _field_stack_stack_num_field_type_22_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'he == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_14_field_type_22_sub_class_id <= _field_stack_stack_num_field_type_22_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'he == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_14_field_type_23_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_23_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'he == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_14_field_type_23_field_type <= _field_stack_stack_num_field_type_23_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'he == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_14_field_type_23_sub_class_id <= _field_stack_stack_num_field_type_23_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'he == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_14_field_type_24_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_24_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'he == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_14_field_type_24_field_type <= _field_stack_stack_num_field_type_24_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'he == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_14_field_type_24_sub_class_id <= _field_stack_stack_num_field_type_24_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'he == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_14_field_type_25_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_25_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'he == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_14_field_type_25_field_type <= _field_stack_stack_num_field_type_25_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'he == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_14_field_type_25_sub_class_id <= _field_stack_stack_num_field_type_25_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'he == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_14_field_type_26_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_26_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'he == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_14_field_type_26_field_type <= _field_stack_stack_num_field_type_26_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'he == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_14_field_type_26_sub_class_id <= _field_stack_stack_num_field_type_26_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'he == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_14_field_type_27_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_27_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'he == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_14_field_type_27_field_type <= _field_stack_stack_num_field_type_27_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'he == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_14_field_type_27_sub_class_id <= _field_stack_stack_num_field_type_27_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'he == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_14_field_type_28_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_28_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'he == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_14_field_type_28_field_type <= _field_stack_stack_num_field_type_28_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'he == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_14_field_type_28_sub_class_id <= _field_stack_stack_num_field_type_28_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'he == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_14_field_type_29_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_29_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'he == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_14_field_type_29_field_type <= _field_stack_stack_num_field_type_29_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'he == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_14_field_type_29_sub_class_id <= _field_stack_stack_num_field_type_29_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'he == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_14_field_type_30_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_30_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'he == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_14_field_type_30_field_type <= _field_stack_stack_num_field_type_30_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'he == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_14_field_type_30_sub_class_id <= _field_stack_stack_num_field_type_30_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'he == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_14_field_type_31_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_31_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'he == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_14_field_type_31_field_type <= _field_stack_stack_num_field_type_31_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'he == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_14_field_type_31_sub_class_id <= _field_stack_stack_num_field_type_31_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'he == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_14_field_type_32_is_repeated <=
              class_meta_rsp_fifo_io_out_bits_class_meta_field_type_32_is_repeated; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'he == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_14_field_type_32_field_type <= _field_stack_stack_num_field_type_32_field_type; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          if (4'he == stack_num) begin // @[Serializerhw.scala 114:45]
            field_stack_14_field_type_32_sub_class_id <= _field_stack_stack_num_field_type_32_sub_class_id; // @[Serializerhw.scala 114:45]
          end
        end
      end
    end
    if (reset) begin // @[Serializerhw.scala 70:28]
      field_num_0 <= 6'h0; // @[Serializerhw.scala 70:28]
    end else if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          field_num_0 <= _GEN_2026;
        end
      end else if (!(_T_8)) begin // @[Conditional.scala 39:67]
        field_num_0 <= _GEN_6502;
      end
    end
    if (reset) begin // @[Serializerhw.scala 70:28]
      field_num_1 <= 6'h0; // @[Serializerhw.scala 70:28]
    end else if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          field_num_1 <= _GEN_2027;
        end
      end else if (!(_T_8)) begin // @[Conditional.scala 39:67]
        field_num_1 <= _GEN_6503;
      end
    end
    if (reset) begin // @[Serializerhw.scala 70:28]
      field_num_2 <= 6'h0; // @[Serializerhw.scala 70:28]
    end else if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          field_num_2 <= _GEN_2028;
        end
      end else if (!(_T_8)) begin // @[Conditional.scala 39:67]
        field_num_2 <= _GEN_6504;
      end
    end
    if (reset) begin // @[Serializerhw.scala 70:28]
      field_num_3 <= 6'h0; // @[Serializerhw.scala 70:28]
    end else if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          field_num_3 <= _GEN_2029;
        end
      end else if (!(_T_8)) begin // @[Conditional.scala 39:67]
        field_num_3 <= _GEN_6505;
      end
    end
    if (reset) begin // @[Serializerhw.scala 70:28]
      field_num_4 <= 6'h0; // @[Serializerhw.scala 70:28]
    end else if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          field_num_4 <= _GEN_2030;
        end
      end else if (!(_T_8)) begin // @[Conditional.scala 39:67]
        field_num_4 <= _GEN_6506;
      end
    end
    if (reset) begin // @[Serializerhw.scala 70:28]
      field_num_5 <= 6'h0; // @[Serializerhw.scala 70:28]
    end else if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          field_num_5 <= _GEN_2031;
        end
      end else if (!(_T_8)) begin // @[Conditional.scala 39:67]
        field_num_5 <= _GEN_6507;
      end
    end
    if (reset) begin // @[Serializerhw.scala 70:28]
      field_num_6 <= 6'h0; // @[Serializerhw.scala 70:28]
    end else if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          field_num_6 <= _GEN_2032;
        end
      end else if (!(_T_8)) begin // @[Conditional.scala 39:67]
        field_num_6 <= _GEN_6508;
      end
    end
    if (reset) begin // @[Serializerhw.scala 70:28]
      field_num_7 <= 6'h0; // @[Serializerhw.scala 70:28]
    end else if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          field_num_7 <= _GEN_2033;
        end
      end else if (!(_T_8)) begin // @[Conditional.scala 39:67]
        field_num_7 <= _GEN_6509;
      end
    end
    if (reset) begin // @[Serializerhw.scala 70:28]
      field_num_8 <= 6'h0; // @[Serializerhw.scala 70:28]
    end else if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          field_num_8 <= _GEN_2034;
        end
      end else if (!(_T_8)) begin // @[Conditional.scala 39:67]
        field_num_8 <= _GEN_6510;
      end
    end
    if (reset) begin // @[Serializerhw.scala 70:28]
      field_num_9 <= 6'h0; // @[Serializerhw.scala 70:28]
    end else if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          field_num_9 <= _GEN_2035;
        end
      end else if (!(_T_8)) begin // @[Conditional.scala 39:67]
        field_num_9 <= _GEN_6511;
      end
    end
    if (reset) begin // @[Serializerhw.scala 70:28]
      field_num_10 <= 6'h0; // @[Serializerhw.scala 70:28]
    end else if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          field_num_10 <= _GEN_2036;
        end
      end else if (!(_T_8)) begin // @[Conditional.scala 39:67]
        field_num_10 <= _GEN_6512;
      end
    end
    if (reset) begin // @[Serializerhw.scala 70:28]
      field_num_11 <= 6'h0; // @[Serializerhw.scala 70:28]
    end else if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          field_num_11 <= _GEN_2037;
        end
      end else if (!(_T_8)) begin // @[Conditional.scala 39:67]
        field_num_11 <= _GEN_6513;
      end
    end
    if (reset) begin // @[Serializerhw.scala 70:28]
      field_num_12 <= 6'h0; // @[Serializerhw.scala 70:28]
    end else if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          field_num_12 <= _GEN_2038;
        end
      end else if (!(_T_8)) begin // @[Conditional.scala 39:67]
        field_num_12 <= _GEN_6514;
      end
    end
    if (reset) begin // @[Serializerhw.scala 70:28]
      field_num_13 <= 6'h0; // @[Serializerhw.scala 70:28]
    end else if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          field_num_13 <= _GEN_2039;
        end
      end else if (!(_T_8)) begin // @[Conditional.scala 39:67]
        field_num_13 <= _GEN_6515;
      end
    end
    if (reset) begin // @[Serializerhw.scala 70:28]
      field_num_14 <= 6'h0; // @[Serializerhw.scala 70:28]
    end else if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          field_num_14 <= _GEN_2040;
        end
      end else if (!(_T_8)) begin // @[Conditional.scala 39:67]
        field_num_14 <= _GEN_6516;
      end
    end
    if (reset) begin // @[Serializerhw.scala 70:28]
      field_num_15 <= 6'h0; // @[Serializerhw.scala 70:28]
    end else if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (_T_6) begin // @[Conditional.scala 39:67]
        if (_T_7) begin // @[Serializerhw.scala 113:52]
          field_num_15 <= _GEN_2041;
        end
      end else if (!(_T_8)) begin // @[Conditional.scala 39:67]
        field_num_15 <= _GEN_6517;
      end
    end
    if (reset) begin // @[Serializerhw.scala 72:33]
      host_base_addr <= 64'h0; // @[Serializerhw.scala 72:33]
    end else if (_T_4) begin // @[Conditional.scala 40:58]
      if (_T_5) begin // @[Serializerhw.scala 102:45]
        host_base_addr <= meta_in_fifo_io_out_bits_host_base_addr; // @[Serializerhw.scala 104:45]
      end
    end else if (_T_6) begin // @[Conditional.scala 39:67]
      if (_T_7) begin // @[Serializerhw.scala 113:52]
        host_base_addr <= _host_base_addr_T_1; // @[Serializerhw.scala 117:45]
      end
    end
    if (reset) begin // @[Serializerhw.scala 73:36]
      current_field_num <= 6'h0; // @[Serializerhw.scala 73:36]
    end else begin
      current_field_num <= _GEN_10631[5:0];
    end
    if (reset) begin // @[Serializerhw.scala 74:33]
      c_sub_metadata_is_repeated <= 1'h0; // @[Serializerhw.scala 74:33]
    end else if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (!(_T_6)) begin // @[Conditional.scala 39:67]
        if (!(_T_8)) begin // @[Conditional.scala 39:67]
          c_sub_metadata_is_repeated <= _GEN_6497;
        end
      end
    end
    if (reset) begin // @[Serializerhw.scala 74:33]
      c_sub_metadata_field_type <= 5'h0; // @[Serializerhw.scala 74:33]
    end else if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (!(_T_6)) begin // @[Conditional.scala 39:67]
        if (!(_T_8)) begin // @[Conditional.scala 39:67]
          c_sub_metadata_field_type <= _GEN_6496;
        end
      end
    end
    if (reset) begin // @[Serializerhw.scala 74:33]
      c_sub_metadata_sub_class_id <= 16'h0; // @[Serializerhw.scala 74:33]
    end else if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (!(_T_6)) begin // @[Conditional.scala 39:67]
        if (!(_T_8)) begin // @[Conditional.scala 39:67]
          c_sub_metadata_sub_class_id <= _GEN_6495;
        end
      end
    end
    if (reset) begin // @[Serializerhw.scala 75:29]
      repeat_num <= 8'h0; // @[Serializerhw.scala 75:29]
    end else begin
      repeat_num <= _GEN_10639[7:0];
    end
    if (reset) begin // @[Serializerhw.scala 76:30]
      stack_num <= 4'h0; // @[Serializerhw.scala 76:30]
    end else if (_T_4) begin // @[Conditional.scala 40:58]
      if (_T_5) begin // @[Serializerhw.scala 102:45]
        stack_num <= 4'h0; // @[Serializerhw.scala 108:45]
      end
    end else if (!(_T_6)) begin // @[Conditional.scala 39:67]
      if (!(_T_8)) begin // @[Conditional.scala 39:67]
        stack_num <= _GEN_6501;
      end
    end
    if (reset) begin // @[Serializerhw.scala 83:38]
      current_field_length <= 32'h0; // @[Serializerhw.scala 83:38]
    end else if (!(_T_4)) begin // @[Conditional.scala 40:58]
      if (!(_T_6)) begin // @[Conditional.scala 39:67]
        if (!(_T_8)) begin // @[Conditional.scala 39:67]
          current_field_length <= _GEN_6518;
        end
      end
    end
    if (reset) begin // @[Serializerhw.scala 86:46]
      state <= 5'h6; // @[Serializerhw.scala 86:46]
    end else if (_T_4) begin // @[Conditional.scala 40:58]
      if (_T_5) begin // @[Serializerhw.scala 102:45]
        state <= 5'h11; // @[Serializerhw.scala 109:45]
      end
    end else if (_T_6) begin // @[Conditional.scala 39:67]
      if (_T_7) begin // @[Serializerhw.scala 113:52]
        state <= 5'h7; // @[Serializerhw.scala 121:45]
      end
    end else if (_T_8) begin // @[Conditional.scala 39:67]
      state <= _GEN_4074;
    end else begin
      state <= _GEN_6492;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  counter = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  counter_1 = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  counter_2 = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  counter_3 = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  field_stack_0_field_type_0_is_repeated = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  field_stack_0_field_type_0_field_type = _RAND_5[4:0];
  _RAND_6 = {1{`RANDOM}};
  field_stack_0_field_type_0_sub_class_id = _RAND_6[15:0];
  _RAND_7 = {1{`RANDOM}};
  field_stack_0_field_type_1_is_repeated = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  field_stack_0_field_type_1_field_type = _RAND_8[4:0];
  _RAND_9 = {1{`RANDOM}};
  field_stack_0_field_type_1_sub_class_id = _RAND_9[15:0];
  _RAND_10 = {1{`RANDOM}};
  field_stack_0_field_type_2_is_repeated = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  field_stack_0_field_type_2_field_type = _RAND_11[4:0];
  _RAND_12 = {1{`RANDOM}};
  field_stack_0_field_type_2_sub_class_id = _RAND_12[15:0];
  _RAND_13 = {1{`RANDOM}};
  field_stack_0_field_type_3_is_repeated = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  field_stack_0_field_type_3_field_type = _RAND_14[4:0];
  _RAND_15 = {1{`RANDOM}};
  field_stack_0_field_type_3_sub_class_id = _RAND_15[15:0];
  _RAND_16 = {1{`RANDOM}};
  field_stack_0_field_type_4_is_repeated = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  field_stack_0_field_type_4_field_type = _RAND_17[4:0];
  _RAND_18 = {1{`RANDOM}};
  field_stack_0_field_type_4_sub_class_id = _RAND_18[15:0];
  _RAND_19 = {1{`RANDOM}};
  field_stack_0_field_type_5_is_repeated = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  field_stack_0_field_type_5_field_type = _RAND_20[4:0];
  _RAND_21 = {1{`RANDOM}};
  field_stack_0_field_type_5_sub_class_id = _RAND_21[15:0];
  _RAND_22 = {1{`RANDOM}};
  field_stack_0_field_type_6_is_repeated = _RAND_22[0:0];
  _RAND_23 = {1{`RANDOM}};
  field_stack_0_field_type_6_field_type = _RAND_23[4:0];
  _RAND_24 = {1{`RANDOM}};
  field_stack_0_field_type_6_sub_class_id = _RAND_24[15:0];
  _RAND_25 = {1{`RANDOM}};
  field_stack_0_field_type_7_is_repeated = _RAND_25[0:0];
  _RAND_26 = {1{`RANDOM}};
  field_stack_0_field_type_7_field_type = _RAND_26[4:0];
  _RAND_27 = {1{`RANDOM}};
  field_stack_0_field_type_7_sub_class_id = _RAND_27[15:0];
  _RAND_28 = {1{`RANDOM}};
  field_stack_0_field_type_8_is_repeated = _RAND_28[0:0];
  _RAND_29 = {1{`RANDOM}};
  field_stack_0_field_type_8_field_type = _RAND_29[4:0];
  _RAND_30 = {1{`RANDOM}};
  field_stack_0_field_type_8_sub_class_id = _RAND_30[15:0];
  _RAND_31 = {1{`RANDOM}};
  field_stack_0_field_type_9_is_repeated = _RAND_31[0:0];
  _RAND_32 = {1{`RANDOM}};
  field_stack_0_field_type_9_field_type = _RAND_32[4:0];
  _RAND_33 = {1{`RANDOM}};
  field_stack_0_field_type_9_sub_class_id = _RAND_33[15:0];
  _RAND_34 = {1{`RANDOM}};
  field_stack_0_field_type_10_is_repeated = _RAND_34[0:0];
  _RAND_35 = {1{`RANDOM}};
  field_stack_0_field_type_10_field_type = _RAND_35[4:0];
  _RAND_36 = {1{`RANDOM}};
  field_stack_0_field_type_10_sub_class_id = _RAND_36[15:0];
  _RAND_37 = {1{`RANDOM}};
  field_stack_0_field_type_11_is_repeated = _RAND_37[0:0];
  _RAND_38 = {1{`RANDOM}};
  field_stack_0_field_type_11_field_type = _RAND_38[4:0];
  _RAND_39 = {1{`RANDOM}};
  field_stack_0_field_type_11_sub_class_id = _RAND_39[15:0];
  _RAND_40 = {1{`RANDOM}};
  field_stack_0_field_type_12_is_repeated = _RAND_40[0:0];
  _RAND_41 = {1{`RANDOM}};
  field_stack_0_field_type_12_field_type = _RAND_41[4:0];
  _RAND_42 = {1{`RANDOM}};
  field_stack_0_field_type_12_sub_class_id = _RAND_42[15:0];
  _RAND_43 = {1{`RANDOM}};
  field_stack_0_field_type_13_is_repeated = _RAND_43[0:0];
  _RAND_44 = {1{`RANDOM}};
  field_stack_0_field_type_13_field_type = _RAND_44[4:0];
  _RAND_45 = {1{`RANDOM}};
  field_stack_0_field_type_13_sub_class_id = _RAND_45[15:0];
  _RAND_46 = {1{`RANDOM}};
  field_stack_0_field_type_14_is_repeated = _RAND_46[0:0];
  _RAND_47 = {1{`RANDOM}};
  field_stack_0_field_type_14_field_type = _RAND_47[4:0];
  _RAND_48 = {1{`RANDOM}};
  field_stack_0_field_type_14_sub_class_id = _RAND_48[15:0];
  _RAND_49 = {1{`RANDOM}};
  field_stack_0_field_type_15_is_repeated = _RAND_49[0:0];
  _RAND_50 = {1{`RANDOM}};
  field_stack_0_field_type_15_field_type = _RAND_50[4:0];
  _RAND_51 = {1{`RANDOM}};
  field_stack_0_field_type_15_sub_class_id = _RAND_51[15:0];
  _RAND_52 = {1{`RANDOM}};
  field_stack_0_field_type_16_is_repeated = _RAND_52[0:0];
  _RAND_53 = {1{`RANDOM}};
  field_stack_0_field_type_16_field_type = _RAND_53[4:0];
  _RAND_54 = {1{`RANDOM}};
  field_stack_0_field_type_16_sub_class_id = _RAND_54[15:0];
  _RAND_55 = {1{`RANDOM}};
  field_stack_0_field_type_17_is_repeated = _RAND_55[0:0];
  _RAND_56 = {1{`RANDOM}};
  field_stack_0_field_type_17_field_type = _RAND_56[4:0];
  _RAND_57 = {1{`RANDOM}};
  field_stack_0_field_type_17_sub_class_id = _RAND_57[15:0];
  _RAND_58 = {1{`RANDOM}};
  field_stack_0_field_type_18_is_repeated = _RAND_58[0:0];
  _RAND_59 = {1{`RANDOM}};
  field_stack_0_field_type_18_field_type = _RAND_59[4:0];
  _RAND_60 = {1{`RANDOM}};
  field_stack_0_field_type_18_sub_class_id = _RAND_60[15:0];
  _RAND_61 = {1{`RANDOM}};
  field_stack_0_field_type_19_is_repeated = _RAND_61[0:0];
  _RAND_62 = {1{`RANDOM}};
  field_stack_0_field_type_19_field_type = _RAND_62[4:0];
  _RAND_63 = {1{`RANDOM}};
  field_stack_0_field_type_19_sub_class_id = _RAND_63[15:0];
  _RAND_64 = {1{`RANDOM}};
  field_stack_0_field_type_20_is_repeated = _RAND_64[0:0];
  _RAND_65 = {1{`RANDOM}};
  field_stack_0_field_type_20_field_type = _RAND_65[4:0];
  _RAND_66 = {1{`RANDOM}};
  field_stack_0_field_type_20_sub_class_id = _RAND_66[15:0];
  _RAND_67 = {1{`RANDOM}};
  field_stack_0_field_type_21_is_repeated = _RAND_67[0:0];
  _RAND_68 = {1{`RANDOM}};
  field_stack_0_field_type_21_field_type = _RAND_68[4:0];
  _RAND_69 = {1{`RANDOM}};
  field_stack_0_field_type_21_sub_class_id = _RAND_69[15:0];
  _RAND_70 = {1{`RANDOM}};
  field_stack_0_field_type_22_is_repeated = _RAND_70[0:0];
  _RAND_71 = {1{`RANDOM}};
  field_stack_0_field_type_22_field_type = _RAND_71[4:0];
  _RAND_72 = {1{`RANDOM}};
  field_stack_0_field_type_22_sub_class_id = _RAND_72[15:0];
  _RAND_73 = {1{`RANDOM}};
  field_stack_0_field_type_23_is_repeated = _RAND_73[0:0];
  _RAND_74 = {1{`RANDOM}};
  field_stack_0_field_type_23_field_type = _RAND_74[4:0];
  _RAND_75 = {1{`RANDOM}};
  field_stack_0_field_type_23_sub_class_id = _RAND_75[15:0];
  _RAND_76 = {1{`RANDOM}};
  field_stack_0_field_type_24_is_repeated = _RAND_76[0:0];
  _RAND_77 = {1{`RANDOM}};
  field_stack_0_field_type_24_field_type = _RAND_77[4:0];
  _RAND_78 = {1{`RANDOM}};
  field_stack_0_field_type_24_sub_class_id = _RAND_78[15:0];
  _RAND_79 = {1{`RANDOM}};
  field_stack_0_field_type_25_is_repeated = _RAND_79[0:0];
  _RAND_80 = {1{`RANDOM}};
  field_stack_0_field_type_25_field_type = _RAND_80[4:0];
  _RAND_81 = {1{`RANDOM}};
  field_stack_0_field_type_25_sub_class_id = _RAND_81[15:0];
  _RAND_82 = {1{`RANDOM}};
  field_stack_0_field_type_26_is_repeated = _RAND_82[0:0];
  _RAND_83 = {1{`RANDOM}};
  field_stack_0_field_type_26_field_type = _RAND_83[4:0];
  _RAND_84 = {1{`RANDOM}};
  field_stack_0_field_type_26_sub_class_id = _RAND_84[15:0];
  _RAND_85 = {1{`RANDOM}};
  field_stack_0_field_type_27_is_repeated = _RAND_85[0:0];
  _RAND_86 = {1{`RANDOM}};
  field_stack_0_field_type_27_field_type = _RAND_86[4:0];
  _RAND_87 = {1{`RANDOM}};
  field_stack_0_field_type_27_sub_class_id = _RAND_87[15:0];
  _RAND_88 = {1{`RANDOM}};
  field_stack_0_field_type_28_is_repeated = _RAND_88[0:0];
  _RAND_89 = {1{`RANDOM}};
  field_stack_0_field_type_28_field_type = _RAND_89[4:0];
  _RAND_90 = {1{`RANDOM}};
  field_stack_0_field_type_28_sub_class_id = _RAND_90[15:0];
  _RAND_91 = {1{`RANDOM}};
  field_stack_0_field_type_29_is_repeated = _RAND_91[0:0];
  _RAND_92 = {1{`RANDOM}};
  field_stack_0_field_type_29_field_type = _RAND_92[4:0];
  _RAND_93 = {1{`RANDOM}};
  field_stack_0_field_type_29_sub_class_id = _RAND_93[15:0];
  _RAND_94 = {1{`RANDOM}};
  field_stack_0_field_type_30_is_repeated = _RAND_94[0:0];
  _RAND_95 = {1{`RANDOM}};
  field_stack_0_field_type_30_field_type = _RAND_95[4:0];
  _RAND_96 = {1{`RANDOM}};
  field_stack_0_field_type_30_sub_class_id = _RAND_96[15:0];
  _RAND_97 = {1{`RANDOM}};
  field_stack_0_field_type_31_is_repeated = _RAND_97[0:0];
  _RAND_98 = {1{`RANDOM}};
  field_stack_0_field_type_31_field_type = _RAND_98[4:0];
  _RAND_99 = {1{`RANDOM}};
  field_stack_0_field_type_31_sub_class_id = _RAND_99[15:0];
  _RAND_100 = {1{`RANDOM}};
  field_stack_0_field_type_32_is_repeated = _RAND_100[0:0];
  _RAND_101 = {1{`RANDOM}};
  field_stack_0_field_type_32_field_type = _RAND_101[4:0];
  _RAND_102 = {1{`RANDOM}};
  field_stack_0_field_type_32_sub_class_id = _RAND_102[15:0];
  _RAND_103 = {1{`RANDOM}};
  field_stack_1_field_type_0_is_repeated = _RAND_103[0:0];
  _RAND_104 = {1{`RANDOM}};
  field_stack_1_field_type_0_field_type = _RAND_104[4:0];
  _RAND_105 = {1{`RANDOM}};
  field_stack_1_field_type_0_sub_class_id = _RAND_105[15:0];
  _RAND_106 = {1{`RANDOM}};
  field_stack_1_field_type_1_is_repeated = _RAND_106[0:0];
  _RAND_107 = {1{`RANDOM}};
  field_stack_1_field_type_1_field_type = _RAND_107[4:0];
  _RAND_108 = {1{`RANDOM}};
  field_stack_1_field_type_1_sub_class_id = _RAND_108[15:0];
  _RAND_109 = {1{`RANDOM}};
  field_stack_1_field_type_2_is_repeated = _RAND_109[0:0];
  _RAND_110 = {1{`RANDOM}};
  field_stack_1_field_type_2_field_type = _RAND_110[4:0];
  _RAND_111 = {1{`RANDOM}};
  field_stack_1_field_type_2_sub_class_id = _RAND_111[15:0];
  _RAND_112 = {1{`RANDOM}};
  field_stack_1_field_type_3_is_repeated = _RAND_112[0:0];
  _RAND_113 = {1{`RANDOM}};
  field_stack_1_field_type_3_field_type = _RAND_113[4:0];
  _RAND_114 = {1{`RANDOM}};
  field_stack_1_field_type_3_sub_class_id = _RAND_114[15:0];
  _RAND_115 = {1{`RANDOM}};
  field_stack_1_field_type_4_is_repeated = _RAND_115[0:0];
  _RAND_116 = {1{`RANDOM}};
  field_stack_1_field_type_4_field_type = _RAND_116[4:0];
  _RAND_117 = {1{`RANDOM}};
  field_stack_1_field_type_4_sub_class_id = _RAND_117[15:0];
  _RAND_118 = {1{`RANDOM}};
  field_stack_1_field_type_5_is_repeated = _RAND_118[0:0];
  _RAND_119 = {1{`RANDOM}};
  field_stack_1_field_type_5_field_type = _RAND_119[4:0];
  _RAND_120 = {1{`RANDOM}};
  field_stack_1_field_type_5_sub_class_id = _RAND_120[15:0];
  _RAND_121 = {1{`RANDOM}};
  field_stack_1_field_type_6_is_repeated = _RAND_121[0:0];
  _RAND_122 = {1{`RANDOM}};
  field_stack_1_field_type_6_field_type = _RAND_122[4:0];
  _RAND_123 = {1{`RANDOM}};
  field_stack_1_field_type_6_sub_class_id = _RAND_123[15:0];
  _RAND_124 = {1{`RANDOM}};
  field_stack_1_field_type_7_is_repeated = _RAND_124[0:0];
  _RAND_125 = {1{`RANDOM}};
  field_stack_1_field_type_7_field_type = _RAND_125[4:0];
  _RAND_126 = {1{`RANDOM}};
  field_stack_1_field_type_7_sub_class_id = _RAND_126[15:0];
  _RAND_127 = {1{`RANDOM}};
  field_stack_1_field_type_8_is_repeated = _RAND_127[0:0];
  _RAND_128 = {1{`RANDOM}};
  field_stack_1_field_type_8_field_type = _RAND_128[4:0];
  _RAND_129 = {1{`RANDOM}};
  field_stack_1_field_type_8_sub_class_id = _RAND_129[15:0];
  _RAND_130 = {1{`RANDOM}};
  field_stack_1_field_type_9_is_repeated = _RAND_130[0:0];
  _RAND_131 = {1{`RANDOM}};
  field_stack_1_field_type_9_field_type = _RAND_131[4:0];
  _RAND_132 = {1{`RANDOM}};
  field_stack_1_field_type_9_sub_class_id = _RAND_132[15:0];
  _RAND_133 = {1{`RANDOM}};
  field_stack_1_field_type_10_is_repeated = _RAND_133[0:0];
  _RAND_134 = {1{`RANDOM}};
  field_stack_1_field_type_10_field_type = _RAND_134[4:0];
  _RAND_135 = {1{`RANDOM}};
  field_stack_1_field_type_10_sub_class_id = _RAND_135[15:0];
  _RAND_136 = {1{`RANDOM}};
  field_stack_1_field_type_11_is_repeated = _RAND_136[0:0];
  _RAND_137 = {1{`RANDOM}};
  field_stack_1_field_type_11_field_type = _RAND_137[4:0];
  _RAND_138 = {1{`RANDOM}};
  field_stack_1_field_type_11_sub_class_id = _RAND_138[15:0];
  _RAND_139 = {1{`RANDOM}};
  field_stack_1_field_type_12_is_repeated = _RAND_139[0:0];
  _RAND_140 = {1{`RANDOM}};
  field_stack_1_field_type_12_field_type = _RAND_140[4:0];
  _RAND_141 = {1{`RANDOM}};
  field_stack_1_field_type_12_sub_class_id = _RAND_141[15:0];
  _RAND_142 = {1{`RANDOM}};
  field_stack_1_field_type_13_is_repeated = _RAND_142[0:0];
  _RAND_143 = {1{`RANDOM}};
  field_stack_1_field_type_13_field_type = _RAND_143[4:0];
  _RAND_144 = {1{`RANDOM}};
  field_stack_1_field_type_13_sub_class_id = _RAND_144[15:0];
  _RAND_145 = {1{`RANDOM}};
  field_stack_1_field_type_14_is_repeated = _RAND_145[0:0];
  _RAND_146 = {1{`RANDOM}};
  field_stack_1_field_type_14_field_type = _RAND_146[4:0];
  _RAND_147 = {1{`RANDOM}};
  field_stack_1_field_type_14_sub_class_id = _RAND_147[15:0];
  _RAND_148 = {1{`RANDOM}};
  field_stack_1_field_type_15_is_repeated = _RAND_148[0:0];
  _RAND_149 = {1{`RANDOM}};
  field_stack_1_field_type_15_field_type = _RAND_149[4:0];
  _RAND_150 = {1{`RANDOM}};
  field_stack_1_field_type_15_sub_class_id = _RAND_150[15:0];
  _RAND_151 = {1{`RANDOM}};
  field_stack_1_field_type_16_is_repeated = _RAND_151[0:0];
  _RAND_152 = {1{`RANDOM}};
  field_stack_1_field_type_16_field_type = _RAND_152[4:0];
  _RAND_153 = {1{`RANDOM}};
  field_stack_1_field_type_16_sub_class_id = _RAND_153[15:0];
  _RAND_154 = {1{`RANDOM}};
  field_stack_1_field_type_17_is_repeated = _RAND_154[0:0];
  _RAND_155 = {1{`RANDOM}};
  field_stack_1_field_type_17_field_type = _RAND_155[4:0];
  _RAND_156 = {1{`RANDOM}};
  field_stack_1_field_type_17_sub_class_id = _RAND_156[15:0];
  _RAND_157 = {1{`RANDOM}};
  field_stack_1_field_type_18_is_repeated = _RAND_157[0:0];
  _RAND_158 = {1{`RANDOM}};
  field_stack_1_field_type_18_field_type = _RAND_158[4:0];
  _RAND_159 = {1{`RANDOM}};
  field_stack_1_field_type_18_sub_class_id = _RAND_159[15:0];
  _RAND_160 = {1{`RANDOM}};
  field_stack_1_field_type_19_is_repeated = _RAND_160[0:0];
  _RAND_161 = {1{`RANDOM}};
  field_stack_1_field_type_19_field_type = _RAND_161[4:0];
  _RAND_162 = {1{`RANDOM}};
  field_stack_1_field_type_19_sub_class_id = _RAND_162[15:0];
  _RAND_163 = {1{`RANDOM}};
  field_stack_1_field_type_20_is_repeated = _RAND_163[0:0];
  _RAND_164 = {1{`RANDOM}};
  field_stack_1_field_type_20_field_type = _RAND_164[4:0];
  _RAND_165 = {1{`RANDOM}};
  field_stack_1_field_type_20_sub_class_id = _RAND_165[15:0];
  _RAND_166 = {1{`RANDOM}};
  field_stack_1_field_type_21_is_repeated = _RAND_166[0:0];
  _RAND_167 = {1{`RANDOM}};
  field_stack_1_field_type_21_field_type = _RAND_167[4:0];
  _RAND_168 = {1{`RANDOM}};
  field_stack_1_field_type_21_sub_class_id = _RAND_168[15:0];
  _RAND_169 = {1{`RANDOM}};
  field_stack_1_field_type_22_is_repeated = _RAND_169[0:0];
  _RAND_170 = {1{`RANDOM}};
  field_stack_1_field_type_22_field_type = _RAND_170[4:0];
  _RAND_171 = {1{`RANDOM}};
  field_stack_1_field_type_22_sub_class_id = _RAND_171[15:0];
  _RAND_172 = {1{`RANDOM}};
  field_stack_1_field_type_23_is_repeated = _RAND_172[0:0];
  _RAND_173 = {1{`RANDOM}};
  field_stack_1_field_type_23_field_type = _RAND_173[4:0];
  _RAND_174 = {1{`RANDOM}};
  field_stack_1_field_type_23_sub_class_id = _RAND_174[15:0];
  _RAND_175 = {1{`RANDOM}};
  field_stack_1_field_type_24_is_repeated = _RAND_175[0:0];
  _RAND_176 = {1{`RANDOM}};
  field_stack_1_field_type_24_field_type = _RAND_176[4:0];
  _RAND_177 = {1{`RANDOM}};
  field_stack_1_field_type_24_sub_class_id = _RAND_177[15:0];
  _RAND_178 = {1{`RANDOM}};
  field_stack_1_field_type_25_is_repeated = _RAND_178[0:0];
  _RAND_179 = {1{`RANDOM}};
  field_stack_1_field_type_25_field_type = _RAND_179[4:0];
  _RAND_180 = {1{`RANDOM}};
  field_stack_1_field_type_25_sub_class_id = _RAND_180[15:0];
  _RAND_181 = {1{`RANDOM}};
  field_stack_1_field_type_26_is_repeated = _RAND_181[0:0];
  _RAND_182 = {1{`RANDOM}};
  field_stack_1_field_type_26_field_type = _RAND_182[4:0];
  _RAND_183 = {1{`RANDOM}};
  field_stack_1_field_type_26_sub_class_id = _RAND_183[15:0];
  _RAND_184 = {1{`RANDOM}};
  field_stack_1_field_type_27_is_repeated = _RAND_184[0:0];
  _RAND_185 = {1{`RANDOM}};
  field_stack_1_field_type_27_field_type = _RAND_185[4:0];
  _RAND_186 = {1{`RANDOM}};
  field_stack_1_field_type_27_sub_class_id = _RAND_186[15:0];
  _RAND_187 = {1{`RANDOM}};
  field_stack_1_field_type_28_is_repeated = _RAND_187[0:0];
  _RAND_188 = {1{`RANDOM}};
  field_stack_1_field_type_28_field_type = _RAND_188[4:0];
  _RAND_189 = {1{`RANDOM}};
  field_stack_1_field_type_28_sub_class_id = _RAND_189[15:0];
  _RAND_190 = {1{`RANDOM}};
  field_stack_1_field_type_29_is_repeated = _RAND_190[0:0];
  _RAND_191 = {1{`RANDOM}};
  field_stack_1_field_type_29_field_type = _RAND_191[4:0];
  _RAND_192 = {1{`RANDOM}};
  field_stack_1_field_type_29_sub_class_id = _RAND_192[15:0];
  _RAND_193 = {1{`RANDOM}};
  field_stack_1_field_type_30_is_repeated = _RAND_193[0:0];
  _RAND_194 = {1{`RANDOM}};
  field_stack_1_field_type_30_field_type = _RAND_194[4:0];
  _RAND_195 = {1{`RANDOM}};
  field_stack_1_field_type_30_sub_class_id = _RAND_195[15:0];
  _RAND_196 = {1{`RANDOM}};
  field_stack_1_field_type_31_is_repeated = _RAND_196[0:0];
  _RAND_197 = {1{`RANDOM}};
  field_stack_1_field_type_31_field_type = _RAND_197[4:0];
  _RAND_198 = {1{`RANDOM}};
  field_stack_1_field_type_31_sub_class_id = _RAND_198[15:0];
  _RAND_199 = {1{`RANDOM}};
  field_stack_1_field_type_32_is_repeated = _RAND_199[0:0];
  _RAND_200 = {1{`RANDOM}};
  field_stack_1_field_type_32_field_type = _RAND_200[4:0];
  _RAND_201 = {1{`RANDOM}};
  field_stack_1_field_type_32_sub_class_id = _RAND_201[15:0];
  _RAND_202 = {1{`RANDOM}};
  field_stack_2_field_type_0_is_repeated = _RAND_202[0:0];
  _RAND_203 = {1{`RANDOM}};
  field_stack_2_field_type_0_field_type = _RAND_203[4:0];
  _RAND_204 = {1{`RANDOM}};
  field_stack_2_field_type_0_sub_class_id = _RAND_204[15:0];
  _RAND_205 = {1{`RANDOM}};
  field_stack_2_field_type_1_is_repeated = _RAND_205[0:0];
  _RAND_206 = {1{`RANDOM}};
  field_stack_2_field_type_1_field_type = _RAND_206[4:0];
  _RAND_207 = {1{`RANDOM}};
  field_stack_2_field_type_1_sub_class_id = _RAND_207[15:0];
  _RAND_208 = {1{`RANDOM}};
  field_stack_2_field_type_2_is_repeated = _RAND_208[0:0];
  _RAND_209 = {1{`RANDOM}};
  field_stack_2_field_type_2_field_type = _RAND_209[4:0];
  _RAND_210 = {1{`RANDOM}};
  field_stack_2_field_type_2_sub_class_id = _RAND_210[15:0];
  _RAND_211 = {1{`RANDOM}};
  field_stack_2_field_type_3_is_repeated = _RAND_211[0:0];
  _RAND_212 = {1{`RANDOM}};
  field_stack_2_field_type_3_field_type = _RAND_212[4:0];
  _RAND_213 = {1{`RANDOM}};
  field_stack_2_field_type_3_sub_class_id = _RAND_213[15:0];
  _RAND_214 = {1{`RANDOM}};
  field_stack_2_field_type_4_is_repeated = _RAND_214[0:0];
  _RAND_215 = {1{`RANDOM}};
  field_stack_2_field_type_4_field_type = _RAND_215[4:0];
  _RAND_216 = {1{`RANDOM}};
  field_stack_2_field_type_4_sub_class_id = _RAND_216[15:0];
  _RAND_217 = {1{`RANDOM}};
  field_stack_2_field_type_5_is_repeated = _RAND_217[0:0];
  _RAND_218 = {1{`RANDOM}};
  field_stack_2_field_type_5_field_type = _RAND_218[4:0];
  _RAND_219 = {1{`RANDOM}};
  field_stack_2_field_type_5_sub_class_id = _RAND_219[15:0];
  _RAND_220 = {1{`RANDOM}};
  field_stack_2_field_type_6_is_repeated = _RAND_220[0:0];
  _RAND_221 = {1{`RANDOM}};
  field_stack_2_field_type_6_field_type = _RAND_221[4:0];
  _RAND_222 = {1{`RANDOM}};
  field_stack_2_field_type_6_sub_class_id = _RAND_222[15:0];
  _RAND_223 = {1{`RANDOM}};
  field_stack_2_field_type_7_is_repeated = _RAND_223[0:0];
  _RAND_224 = {1{`RANDOM}};
  field_stack_2_field_type_7_field_type = _RAND_224[4:0];
  _RAND_225 = {1{`RANDOM}};
  field_stack_2_field_type_7_sub_class_id = _RAND_225[15:0];
  _RAND_226 = {1{`RANDOM}};
  field_stack_2_field_type_8_is_repeated = _RAND_226[0:0];
  _RAND_227 = {1{`RANDOM}};
  field_stack_2_field_type_8_field_type = _RAND_227[4:0];
  _RAND_228 = {1{`RANDOM}};
  field_stack_2_field_type_8_sub_class_id = _RAND_228[15:0];
  _RAND_229 = {1{`RANDOM}};
  field_stack_2_field_type_9_is_repeated = _RAND_229[0:0];
  _RAND_230 = {1{`RANDOM}};
  field_stack_2_field_type_9_field_type = _RAND_230[4:0];
  _RAND_231 = {1{`RANDOM}};
  field_stack_2_field_type_9_sub_class_id = _RAND_231[15:0];
  _RAND_232 = {1{`RANDOM}};
  field_stack_2_field_type_10_is_repeated = _RAND_232[0:0];
  _RAND_233 = {1{`RANDOM}};
  field_stack_2_field_type_10_field_type = _RAND_233[4:0];
  _RAND_234 = {1{`RANDOM}};
  field_stack_2_field_type_10_sub_class_id = _RAND_234[15:0];
  _RAND_235 = {1{`RANDOM}};
  field_stack_2_field_type_11_is_repeated = _RAND_235[0:0];
  _RAND_236 = {1{`RANDOM}};
  field_stack_2_field_type_11_field_type = _RAND_236[4:0];
  _RAND_237 = {1{`RANDOM}};
  field_stack_2_field_type_11_sub_class_id = _RAND_237[15:0];
  _RAND_238 = {1{`RANDOM}};
  field_stack_2_field_type_12_is_repeated = _RAND_238[0:0];
  _RAND_239 = {1{`RANDOM}};
  field_stack_2_field_type_12_field_type = _RAND_239[4:0];
  _RAND_240 = {1{`RANDOM}};
  field_stack_2_field_type_12_sub_class_id = _RAND_240[15:0];
  _RAND_241 = {1{`RANDOM}};
  field_stack_2_field_type_13_is_repeated = _RAND_241[0:0];
  _RAND_242 = {1{`RANDOM}};
  field_stack_2_field_type_13_field_type = _RAND_242[4:0];
  _RAND_243 = {1{`RANDOM}};
  field_stack_2_field_type_13_sub_class_id = _RAND_243[15:0];
  _RAND_244 = {1{`RANDOM}};
  field_stack_2_field_type_14_is_repeated = _RAND_244[0:0];
  _RAND_245 = {1{`RANDOM}};
  field_stack_2_field_type_14_field_type = _RAND_245[4:0];
  _RAND_246 = {1{`RANDOM}};
  field_stack_2_field_type_14_sub_class_id = _RAND_246[15:0];
  _RAND_247 = {1{`RANDOM}};
  field_stack_2_field_type_15_is_repeated = _RAND_247[0:0];
  _RAND_248 = {1{`RANDOM}};
  field_stack_2_field_type_15_field_type = _RAND_248[4:0];
  _RAND_249 = {1{`RANDOM}};
  field_stack_2_field_type_15_sub_class_id = _RAND_249[15:0];
  _RAND_250 = {1{`RANDOM}};
  field_stack_2_field_type_16_is_repeated = _RAND_250[0:0];
  _RAND_251 = {1{`RANDOM}};
  field_stack_2_field_type_16_field_type = _RAND_251[4:0];
  _RAND_252 = {1{`RANDOM}};
  field_stack_2_field_type_16_sub_class_id = _RAND_252[15:0];
  _RAND_253 = {1{`RANDOM}};
  field_stack_2_field_type_17_is_repeated = _RAND_253[0:0];
  _RAND_254 = {1{`RANDOM}};
  field_stack_2_field_type_17_field_type = _RAND_254[4:0];
  _RAND_255 = {1{`RANDOM}};
  field_stack_2_field_type_17_sub_class_id = _RAND_255[15:0];
  _RAND_256 = {1{`RANDOM}};
  field_stack_2_field_type_18_is_repeated = _RAND_256[0:0];
  _RAND_257 = {1{`RANDOM}};
  field_stack_2_field_type_18_field_type = _RAND_257[4:0];
  _RAND_258 = {1{`RANDOM}};
  field_stack_2_field_type_18_sub_class_id = _RAND_258[15:0];
  _RAND_259 = {1{`RANDOM}};
  field_stack_2_field_type_19_is_repeated = _RAND_259[0:0];
  _RAND_260 = {1{`RANDOM}};
  field_stack_2_field_type_19_field_type = _RAND_260[4:0];
  _RAND_261 = {1{`RANDOM}};
  field_stack_2_field_type_19_sub_class_id = _RAND_261[15:0];
  _RAND_262 = {1{`RANDOM}};
  field_stack_2_field_type_20_is_repeated = _RAND_262[0:0];
  _RAND_263 = {1{`RANDOM}};
  field_stack_2_field_type_20_field_type = _RAND_263[4:0];
  _RAND_264 = {1{`RANDOM}};
  field_stack_2_field_type_20_sub_class_id = _RAND_264[15:0];
  _RAND_265 = {1{`RANDOM}};
  field_stack_2_field_type_21_is_repeated = _RAND_265[0:0];
  _RAND_266 = {1{`RANDOM}};
  field_stack_2_field_type_21_field_type = _RAND_266[4:0];
  _RAND_267 = {1{`RANDOM}};
  field_stack_2_field_type_21_sub_class_id = _RAND_267[15:0];
  _RAND_268 = {1{`RANDOM}};
  field_stack_2_field_type_22_is_repeated = _RAND_268[0:0];
  _RAND_269 = {1{`RANDOM}};
  field_stack_2_field_type_22_field_type = _RAND_269[4:0];
  _RAND_270 = {1{`RANDOM}};
  field_stack_2_field_type_22_sub_class_id = _RAND_270[15:0];
  _RAND_271 = {1{`RANDOM}};
  field_stack_2_field_type_23_is_repeated = _RAND_271[0:0];
  _RAND_272 = {1{`RANDOM}};
  field_stack_2_field_type_23_field_type = _RAND_272[4:0];
  _RAND_273 = {1{`RANDOM}};
  field_stack_2_field_type_23_sub_class_id = _RAND_273[15:0];
  _RAND_274 = {1{`RANDOM}};
  field_stack_2_field_type_24_is_repeated = _RAND_274[0:0];
  _RAND_275 = {1{`RANDOM}};
  field_stack_2_field_type_24_field_type = _RAND_275[4:0];
  _RAND_276 = {1{`RANDOM}};
  field_stack_2_field_type_24_sub_class_id = _RAND_276[15:0];
  _RAND_277 = {1{`RANDOM}};
  field_stack_2_field_type_25_is_repeated = _RAND_277[0:0];
  _RAND_278 = {1{`RANDOM}};
  field_stack_2_field_type_25_field_type = _RAND_278[4:0];
  _RAND_279 = {1{`RANDOM}};
  field_stack_2_field_type_25_sub_class_id = _RAND_279[15:0];
  _RAND_280 = {1{`RANDOM}};
  field_stack_2_field_type_26_is_repeated = _RAND_280[0:0];
  _RAND_281 = {1{`RANDOM}};
  field_stack_2_field_type_26_field_type = _RAND_281[4:0];
  _RAND_282 = {1{`RANDOM}};
  field_stack_2_field_type_26_sub_class_id = _RAND_282[15:0];
  _RAND_283 = {1{`RANDOM}};
  field_stack_2_field_type_27_is_repeated = _RAND_283[0:0];
  _RAND_284 = {1{`RANDOM}};
  field_stack_2_field_type_27_field_type = _RAND_284[4:0];
  _RAND_285 = {1{`RANDOM}};
  field_stack_2_field_type_27_sub_class_id = _RAND_285[15:0];
  _RAND_286 = {1{`RANDOM}};
  field_stack_2_field_type_28_is_repeated = _RAND_286[0:0];
  _RAND_287 = {1{`RANDOM}};
  field_stack_2_field_type_28_field_type = _RAND_287[4:0];
  _RAND_288 = {1{`RANDOM}};
  field_stack_2_field_type_28_sub_class_id = _RAND_288[15:0];
  _RAND_289 = {1{`RANDOM}};
  field_stack_2_field_type_29_is_repeated = _RAND_289[0:0];
  _RAND_290 = {1{`RANDOM}};
  field_stack_2_field_type_29_field_type = _RAND_290[4:0];
  _RAND_291 = {1{`RANDOM}};
  field_stack_2_field_type_29_sub_class_id = _RAND_291[15:0];
  _RAND_292 = {1{`RANDOM}};
  field_stack_2_field_type_30_is_repeated = _RAND_292[0:0];
  _RAND_293 = {1{`RANDOM}};
  field_stack_2_field_type_30_field_type = _RAND_293[4:0];
  _RAND_294 = {1{`RANDOM}};
  field_stack_2_field_type_30_sub_class_id = _RAND_294[15:0];
  _RAND_295 = {1{`RANDOM}};
  field_stack_2_field_type_31_is_repeated = _RAND_295[0:0];
  _RAND_296 = {1{`RANDOM}};
  field_stack_2_field_type_31_field_type = _RAND_296[4:0];
  _RAND_297 = {1{`RANDOM}};
  field_stack_2_field_type_31_sub_class_id = _RAND_297[15:0];
  _RAND_298 = {1{`RANDOM}};
  field_stack_2_field_type_32_is_repeated = _RAND_298[0:0];
  _RAND_299 = {1{`RANDOM}};
  field_stack_2_field_type_32_field_type = _RAND_299[4:0];
  _RAND_300 = {1{`RANDOM}};
  field_stack_2_field_type_32_sub_class_id = _RAND_300[15:0];
  _RAND_301 = {1{`RANDOM}};
  field_stack_3_field_type_0_is_repeated = _RAND_301[0:0];
  _RAND_302 = {1{`RANDOM}};
  field_stack_3_field_type_0_field_type = _RAND_302[4:0];
  _RAND_303 = {1{`RANDOM}};
  field_stack_3_field_type_0_sub_class_id = _RAND_303[15:0];
  _RAND_304 = {1{`RANDOM}};
  field_stack_3_field_type_1_is_repeated = _RAND_304[0:0];
  _RAND_305 = {1{`RANDOM}};
  field_stack_3_field_type_1_field_type = _RAND_305[4:0];
  _RAND_306 = {1{`RANDOM}};
  field_stack_3_field_type_1_sub_class_id = _RAND_306[15:0];
  _RAND_307 = {1{`RANDOM}};
  field_stack_3_field_type_2_is_repeated = _RAND_307[0:0];
  _RAND_308 = {1{`RANDOM}};
  field_stack_3_field_type_2_field_type = _RAND_308[4:0];
  _RAND_309 = {1{`RANDOM}};
  field_stack_3_field_type_2_sub_class_id = _RAND_309[15:0];
  _RAND_310 = {1{`RANDOM}};
  field_stack_3_field_type_3_is_repeated = _RAND_310[0:0];
  _RAND_311 = {1{`RANDOM}};
  field_stack_3_field_type_3_field_type = _RAND_311[4:0];
  _RAND_312 = {1{`RANDOM}};
  field_stack_3_field_type_3_sub_class_id = _RAND_312[15:0];
  _RAND_313 = {1{`RANDOM}};
  field_stack_3_field_type_4_is_repeated = _RAND_313[0:0];
  _RAND_314 = {1{`RANDOM}};
  field_stack_3_field_type_4_field_type = _RAND_314[4:0];
  _RAND_315 = {1{`RANDOM}};
  field_stack_3_field_type_4_sub_class_id = _RAND_315[15:0];
  _RAND_316 = {1{`RANDOM}};
  field_stack_3_field_type_5_is_repeated = _RAND_316[0:0];
  _RAND_317 = {1{`RANDOM}};
  field_stack_3_field_type_5_field_type = _RAND_317[4:0];
  _RAND_318 = {1{`RANDOM}};
  field_stack_3_field_type_5_sub_class_id = _RAND_318[15:0];
  _RAND_319 = {1{`RANDOM}};
  field_stack_3_field_type_6_is_repeated = _RAND_319[0:0];
  _RAND_320 = {1{`RANDOM}};
  field_stack_3_field_type_6_field_type = _RAND_320[4:0];
  _RAND_321 = {1{`RANDOM}};
  field_stack_3_field_type_6_sub_class_id = _RAND_321[15:0];
  _RAND_322 = {1{`RANDOM}};
  field_stack_3_field_type_7_is_repeated = _RAND_322[0:0];
  _RAND_323 = {1{`RANDOM}};
  field_stack_3_field_type_7_field_type = _RAND_323[4:0];
  _RAND_324 = {1{`RANDOM}};
  field_stack_3_field_type_7_sub_class_id = _RAND_324[15:0];
  _RAND_325 = {1{`RANDOM}};
  field_stack_3_field_type_8_is_repeated = _RAND_325[0:0];
  _RAND_326 = {1{`RANDOM}};
  field_stack_3_field_type_8_field_type = _RAND_326[4:0];
  _RAND_327 = {1{`RANDOM}};
  field_stack_3_field_type_8_sub_class_id = _RAND_327[15:0];
  _RAND_328 = {1{`RANDOM}};
  field_stack_3_field_type_9_is_repeated = _RAND_328[0:0];
  _RAND_329 = {1{`RANDOM}};
  field_stack_3_field_type_9_field_type = _RAND_329[4:0];
  _RAND_330 = {1{`RANDOM}};
  field_stack_3_field_type_9_sub_class_id = _RAND_330[15:0];
  _RAND_331 = {1{`RANDOM}};
  field_stack_3_field_type_10_is_repeated = _RAND_331[0:0];
  _RAND_332 = {1{`RANDOM}};
  field_stack_3_field_type_10_field_type = _RAND_332[4:0];
  _RAND_333 = {1{`RANDOM}};
  field_stack_3_field_type_10_sub_class_id = _RAND_333[15:0];
  _RAND_334 = {1{`RANDOM}};
  field_stack_3_field_type_11_is_repeated = _RAND_334[0:0];
  _RAND_335 = {1{`RANDOM}};
  field_stack_3_field_type_11_field_type = _RAND_335[4:0];
  _RAND_336 = {1{`RANDOM}};
  field_stack_3_field_type_11_sub_class_id = _RAND_336[15:0];
  _RAND_337 = {1{`RANDOM}};
  field_stack_3_field_type_12_is_repeated = _RAND_337[0:0];
  _RAND_338 = {1{`RANDOM}};
  field_stack_3_field_type_12_field_type = _RAND_338[4:0];
  _RAND_339 = {1{`RANDOM}};
  field_stack_3_field_type_12_sub_class_id = _RAND_339[15:0];
  _RAND_340 = {1{`RANDOM}};
  field_stack_3_field_type_13_is_repeated = _RAND_340[0:0];
  _RAND_341 = {1{`RANDOM}};
  field_stack_3_field_type_13_field_type = _RAND_341[4:0];
  _RAND_342 = {1{`RANDOM}};
  field_stack_3_field_type_13_sub_class_id = _RAND_342[15:0];
  _RAND_343 = {1{`RANDOM}};
  field_stack_3_field_type_14_is_repeated = _RAND_343[0:0];
  _RAND_344 = {1{`RANDOM}};
  field_stack_3_field_type_14_field_type = _RAND_344[4:0];
  _RAND_345 = {1{`RANDOM}};
  field_stack_3_field_type_14_sub_class_id = _RAND_345[15:0];
  _RAND_346 = {1{`RANDOM}};
  field_stack_3_field_type_15_is_repeated = _RAND_346[0:0];
  _RAND_347 = {1{`RANDOM}};
  field_stack_3_field_type_15_field_type = _RAND_347[4:0];
  _RAND_348 = {1{`RANDOM}};
  field_stack_3_field_type_15_sub_class_id = _RAND_348[15:0];
  _RAND_349 = {1{`RANDOM}};
  field_stack_3_field_type_16_is_repeated = _RAND_349[0:0];
  _RAND_350 = {1{`RANDOM}};
  field_stack_3_field_type_16_field_type = _RAND_350[4:0];
  _RAND_351 = {1{`RANDOM}};
  field_stack_3_field_type_16_sub_class_id = _RAND_351[15:0];
  _RAND_352 = {1{`RANDOM}};
  field_stack_3_field_type_17_is_repeated = _RAND_352[0:0];
  _RAND_353 = {1{`RANDOM}};
  field_stack_3_field_type_17_field_type = _RAND_353[4:0];
  _RAND_354 = {1{`RANDOM}};
  field_stack_3_field_type_17_sub_class_id = _RAND_354[15:0];
  _RAND_355 = {1{`RANDOM}};
  field_stack_3_field_type_18_is_repeated = _RAND_355[0:0];
  _RAND_356 = {1{`RANDOM}};
  field_stack_3_field_type_18_field_type = _RAND_356[4:0];
  _RAND_357 = {1{`RANDOM}};
  field_stack_3_field_type_18_sub_class_id = _RAND_357[15:0];
  _RAND_358 = {1{`RANDOM}};
  field_stack_3_field_type_19_is_repeated = _RAND_358[0:0];
  _RAND_359 = {1{`RANDOM}};
  field_stack_3_field_type_19_field_type = _RAND_359[4:0];
  _RAND_360 = {1{`RANDOM}};
  field_stack_3_field_type_19_sub_class_id = _RAND_360[15:0];
  _RAND_361 = {1{`RANDOM}};
  field_stack_3_field_type_20_is_repeated = _RAND_361[0:0];
  _RAND_362 = {1{`RANDOM}};
  field_stack_3_field_type_20_field_type = _RAND_362[4:0];
  _RAND_363 = {1{`RANDOM}};
  field_stack_3_field_type_20_sub_class_id = _RAND_363[15:0];
  _RAND_364 = {1{`RANDOM}};
  field_stack_3_field_type_21_is_repeated = _RAND_364[0:0];
  _RAND_365 = {1{`RANDOM}};
  field_stack_3_field_type_21_field_type = _RAND_365[4:0];
  _RAND_366 = {1{`RANDOM}};
  field_stack_3_field_type_21_sub_class_id = _RAND_366[15:0];
  _RAND_367 = {1{`RANDOM}};
  field_stack_3_field_type_22_is_repeated = _RAND_367[0:0];
  _RAND_368 = {1{`RANDOM}};
  field_stack_3_field_type_22_field_type = _RAND_368[4:0];
  _RAND_369 = {1{`RANDOM}};
  field_stack_3_field_type_22_sub_class_id = _RAND_369[15:0];
  _RAND_370 = {1{`RANDOM}};
  field_stack_3_field_type_23_is_repeated = _RAND_370[0:0];
  _RAND_371 = {1{`RANDOM}};
  field_stack_3_field_type_23_field_type = _RAND_371[4:0];
  _RAND_372 = {1{`RANDOM}};
  field_stack_3_field_type_23_sub_class_id = _RAND_372[15:0];
  _RAND_373 = {1{`RANDOM}};
  field_stack_3_field_type_24_is_repeated = _RAND_373[0:0];
  _RAND_374 = {1{`RANDOM}};
  field_stack_3_field_type_24_field_type = _RAND_374[4:0];
  _RAND_375 = {1{`RANDOM}};
  field_stack_3_field_type_24_sub_class_id = _RAND_375[15:0];
  _RAND_376 = {1{`RANDOM}};
  field_stack_3_field_type_25_is_repeated = _RAND_376[0:0];
  _RAND_377 = {1{`RANDOM}};
  field_stack_3_field_type_25_field_type = _RAND_377[4:0];
  _RAND_378 = {1{`RANDOM}};
  field_stack_3_field_type_25_sub_class_id = _RAND_378[15:0];
  _RAND_379 = {1{`RANDOM}};
  field_stack_3_field_type_26_is_repeated = _RAND_379[0:0];
  _RAND_380 = {1{`RANDOM}};
  field_stack_3_field_type_26_field_type = _RAND_380[4:0];
  _RAND_381 = {1{`RANDOM}};
  field_stack_3_field_type_26_sub_class_id = _RAND_381[15:0];
  _RAND_382 = {1{`RANDOM}};
  field_stack_3_field_type_27_is_repeated = _RAND_382[0:0];
  _RAND_383 = {1{`RANDOM}};
  field_stack_3_field_type_27_field_type = _RAND_383[4:0];
  _RAND_384 = {1{`RANDOM}};
  field_stack_3_field_type_27_sub_class_id = _RAND_384[15:0];
  _RAND_385 = {1{`RANDOM}};
  field_stack_3_field_type_28_is_repeated = _RAND_385[0:0];
  _RAND_386 = {1{`RANDOM}};
  field_stack_3_field_type_28_field_type = _RAND_386[4:0];
  _RAND_387 = {1{`RANDOM}};
  field_stack_3_field_type_28_sub_class_id = _RAND_387[15:0];
  _RAND_388 = {1{`RANDOM}};
  field_stack_3_field_type_29_is_repeated = _RAND_388[0:0];
  _RAND_389 = {1{`RANDOM}};
  field_stack_3_field_type_29_field_type = _RAND_389[4:0];
  _RAND_390 = {1{`RANDOM}};
  field_stack_3_field_type_29_sub_class_id = _RAND_390[15:0];
  _RAND_391 = {1{`RANDOM}};
  field_stack_3_field_type_30_is_repeated = _RAND_391[0:0];
  _RAND_392 = {1{`RANDOM}};
  field_stack_3_field_type_30_field_type = _RAND_392[4:0];
  _RAND_393 = {1{`RANDOM}};
  field_stack_3_field_type_30_sub_class_id = _RAND_393[15:0];
  _RAND_394 = {1{`RANDOM}};
  field_stack_3_field_type_31_is_repeated = _RAND_394[0:0];
  _RAND_395 = {1{`RANDOM}};
  field_stack_3_field_type_31_field_type = _RAND_395[4:0];
  _RAND_396 = {1{`RANDOM}};
  field_stack_3_field_type_31_sub_class_id = _RAND_396[15:0];
  _RAND_397 = {1{`RANDOM}};
  field_stack_3_field_type_32_is_repeated = _RAND_397[0:0];
  _RAND_398 = {1{`RANDOM}};
  field_stack_3_field_type_32_field_type = _RAND_398[4:0];
  _RAND_399 = {1{`RANDOM}};
  field_stack_3_field_type_32_sub_class_id = _RAND_399[15:0];
  _RAND_400 = {1{`RANDOM}};
  field_stack_4_field_type_0_is_repeated = _RAND_400[0:0];
  _RAND_401 = {1{`RANDOM}};
  field_stack_4_field_type_0_field_type = _RAND_401[4:0];
  _RAND_402 = {1{`RANDOM}};
  field_stack_4_field_type_0_sub_class_id = _RAND_402[15:0];
  _RAND_403 = {1{`RANDOM}};
  field_stack_4_field_type_1_is_repeated = _RAND_403[0:0];
  _RAND_404 = {1{`RANDOM}};
  field_stack_4_field_type_1_field_type = _RAND_404[4:0];
  _RAND_405 = {1{`RANDOM}};
  field_stack_4_field_type_1_sub_class_id = _RAND_405[15:0];
  _RAND_406 = {1{`RANDOM}};
  field_stack_4_field_type_2_is_repeated = _RAND_406[0:0];
  _RAND_407 = {1{`RANDOM}};
  field_stack_4_field_type_2_field_type = _RAND_407[4:0];
  _RAND_408 = {1{`RANDOM}};
  field_stack_4_field_type_2_sub_class_id = _RAND_408[15:0];
  _RAND_409 = {1{`RANDOM}};
  field_stack_4_field_type_3_is_repeated = _RAND_409[0:0];
  _RAND_410 = {1{`RANDOM}};
  field_stack_4_field_type_3_field_type = _RAND_410[4:0];
  _RAND_411 = {1{`RANDOM}};
  field_stack_4_field_type_3_sub_class_id = _RAND_411[15:0];
  _RAND_412 = {1{`RANDOM}};
  field_stack_4_field_type_4_is_repeated = _RAND_412[0:0];
  _RAND_413 = {1{`RANDOM}};
  field_stack_4_field_type_4_field_type = _RAND_413[4:0];
  _RAND_414 = {1{`RANDOM}};
  field_stack_4_field_type_4_sub_class_id = _RAND_414[15:0];
  _RAND_415 = {1{`RANDOM}};
  field_stack_4_field_type_5_is_repeated = _RAND_415[0:0];
  _RAND_416 = {1{`RANDOM}};
  field_stack_4_field_type_5_field_type = _RAND_416[4:0];
  _RAND_417 = {1{`RANDOM}};
  field_stack_4_field_type_5_sub_class_id = _RAND_417[15:0];
  _RAND_418 = {1{`RANDOM}};
  field_stack_4_field_type_6_is_repeated = _RAND_418[0:0];
  _RAND_419 = {1{`RANDOM}};
  field_stack_4_field_type_6_field_type = _RAND_419[4:0];
  _RAND_420 = {1{`RANDOM}};
  field_stack_4_field_type_6_sub_class_id = _RAND_420[15:0];
  _RAND_421 = {1{`RANDOM}};
  field_stack_4_field_type_7_is_repeated = _RAND_421[0:0];
  _RAND_422 = {1{`RANDOM}};
  field_stack_4_field_type_7_field_type = _RAND_422[4:0];
  _RAND_423 = {1{`RANDOM}};
  field_stack_4_field_type_7_sub_class_id = _RAND_423[15:0];
  _RAND_424 = {1{`RANDOM}};
  field_stack_4_field_type_8_is_repeated = _RAND_424[0:0];
  _RAND_425 = {1{`RANDOM}};
  field_stack_4_field_type_8_field_type = _RAND_425[4:0];
  _RAND_426 = {1{`RANDOM}};
  field_stack_4_field_type_8_sub_class_id = _RAND_426[15:0];
  _RAND_427 = {1{`RANDOM}};
  field_stack_4_field_type_9_is_repeated = _RAND_427[0:0];
  _RAND_428 = {1{`RANDOM}};
  field_stack_4_field_type_9_field_type = _RAND_428[4:0];
  _RAND_429 = {1{`RANDOM}};
  field_stack_4_field_type_9_sub_class_id = _RAND_429[15:0];
  _RAND_430 = {1{`RANDOM}};
  field_stack_4_field_type_10_is_repeated = _RAND_430[0:0];
  _RAND_431 = {1{`RANDOM}};
  field_stack_4_field_type_10_field_type = _RAND_431[4:0];
  _RAND_432 = {1{`RANDOM}};
  field_stack_4_field_type_10_sub_class_id = _RAND_432[15:0];
  _RAND_433 = {1{`RANDOM}};
  field_stack_4_field_type_11_is_repeated = _RAND_433[0:0];
  _RAND_434 = {1{`RANDOM}};
  field_stack_4_field_type_11_field_type = _RAND_434[4:0];
  _RAND_435 = {1{`RANDOM}};
  field_stack_4_field_type_11_sub_class_id = _RAND_435[15:0];
  _RAND_436 = {1{`RANDOM}};
  field_stack_4_field_type_12_is_repeated = _RAND_436[0:0];
  _RAND_437 = {1{`RANDOM}};
  field_stack_4_field_type_12_field_type = _RAND_437[4:0];
  _RAND_438 = {1{`RANDOM}};
  field_stack_4_field_type_12_sub_class_id = _RAND_438[15:0];
  _RAND_439 = {1{`RANDOM}};
  field_stack_4_field_type_13_is_repeated = _RAND_439[0:0];
  _RAND_440 = {1{`RANDOM}};
  field_stack_4_field_type_13_field_type = _RAND_440[4:0];
  _RAND_441 = {1{`RANDOM}};
  field_stack_4_field_type_13_sub_class_id = _RAND_441[15:0];
  _RAND_442 = {1{`RANDOM}};
  field_stack_4_field_type_14_is_repeated = _RAND_442[0:0];
  _RAND_443 = {1{`RANDOM}};
  field_stack_4_field_type_14_field_type = _RAND_443[4:0];
  _RAND_444 = {1{`RANDOM}};
  field_stack_4_field_type_14_sub_class_id = _RAND_444[15:0];
  _RAND_445 = {1{`RANDOM}};
  field_stack_4_field_type_15_is_repeated = _RAND_445[0:0];
  _RAND_446 = {1{`RANDOM}};
  field_stack_4_field_type_15_field_type = _RAND_446[4:0];
  _RAND_447 = {1{`RANDOM}};
  field_stack_4_field_type_15_sub_class_id = _RAND_447[15:0];
  _RAND_448 = {1{`RANDOM}};
  field_stack_4_field_type_16_is_repeated = _RAND_448[0:0];
  _RAND_449 = {1{`RANDOM}};
  field_stack_4_field_type_16_field_type = _RAND_449[4:0];
  _RAND_450 = {1{`RANDOM}};
  field_stack_4_field_type_16_sub_class_id = _RAND_450[15:0];
  _RAND_451 = {1{`RANDOM}};
  field_stack_4_field_type_17_is_repeated = _RAND_451[0:0];
  _RAND_452 = {1{`RANDOM}};
  field_stack_4_field_type_17_field_type = _RAND_452[4:0];
  _RAND_453 = {1{`RANDOM}};
  field_stack_4_field_type_17_sub_class_id = _RAND_453[15:0];
  _RAND_454 = {1{`RANDOM}};
  field_stack_4_field_type_18_is_repeated = _RAND_454[0:0];
  _RAND_455 = {1{`RANDOM}};
  field_stack_4_field_type_18_field_type = _RAND_455[4:0];
  _RAND_456 = {1{`RANDOM}};
  field_stack_4_field_type_18_sub_class_id = _RAND_456[15:0];
  _RAND_457 = {1{`RANDOM}};
  field_stack_4_field_type_19_is_repeated = _RAND_457[0:0];
  _RAND_458 = {1{`RANDOM}};
  field_stack_4_field_type_19_field_type = _RAND_458[4:0];
  _RAND_459 = {1{`RANDOM}};
  field_stack_4_field_type_19_sub_class_id = _RAND_459[15:0];
  _RAND_460 = {1{`RANDOM}};
  field_stack_4_field_type_20_is_repeated = _RAND_460[0:0];
  _RAND_461 = {1{`RANDOM}};
  field_stack_4_field_type_20_field_type = _RAND_461[4:0];
  _RAND_462 = {1{`RANDOM}};
  field_stack_4_field_type_20_sub_class_id = _RAND_462[15:0];
  _RAND_463 = {1{`RANDOM}};
  field_stack_4_field_type_21_is_repeated = _RAND_463[0:0];
  _RAND_464 = {1{`RANDOM}};
  field_stack_4_field_type_21_field_type = _RAND_464[4:0];
  _RAND_465 = {1{`RANDOM}};
  field_stack_4_field_type_21_sub_class_id = _RAND_465[15:0];
  _RAND_466 = {1{`RANDOM}};
  field_stack_4_field_type_22_is_repeated = _RAND_466[0:0];
  _RAND_467 = {1{`RANDOM}};
  field_stack_4_field_type_22_field_type = _RAND_467[4:0];
  _RAND_468 = {1{`RANDOM}};
  field_stack_4_field_type_22_sub_class_id = _RAND_468[15:0];
  _RAND_469 = {1{`RANDOM}};
  field_stack_4_field_type_23_is_repeated = _RAND_469[0:0];
  _RAND_470 = {1{`RANDOM}};
  field_stack_4_field_type_23_field_type = _RAND_470[4:0];
  _RAND_471 = {1{`RANDOM}};
  field_stack_4_field_type_23_sub_class_id = _RAND_471[15:0];
  _RAND_472 = {1{`RANDOM}};
  field_stack_4_field_type_24_is_repeated = _RAND_472[0:0];
  _RAND_473 = {1{`RANDOM}};
  field_stack_4_field_type_24_field_type = _RAND_473[4:0];
  _RAND_474 = {1{`RANDOM}};
  field_stack_4_field_type_24_sub_class_id = _RAND_474[15:0];
  _RAND_475 = {1{`RANDOM}};
  field_stack_4_field_type_25_is_repeated = _RAND_475[0:0];
  _RAND_476 = {1{`RANDOM}};
  field_stack_4_field_type_25_field_type = _RAND_476[4:0];
  _RAND_477 = {1{`RANDOM}};
  field_stack_4_field_type_25_sub_class_id = _RAND_477[15:0];
  _RAND_478 = {1{`RANDOM}};
  field_stack_4_field_type_26_is_repeated = _RAND_478[0:0];
  _RAND_479 = {1{`RANDOM}};
  field_stack_4_field_type_26_field_type = _RAND_479[4:0];
  _RAND_480 = {1{`RANDOM}};
  field_stack_4_field_type_26_sub_class_id = _RAND_480[15:0];
  _RAND_481 = {1{`RANDOM}};
  field_stack_4_field_type_27_is_repeated = _RAND_481[0:0];
  _RAND_482 = {1{`RANDOM}};
  field_stack_4_field_type_27_field_type = _RAND_482[4:0];
  _RAND_483 = {1{`RANDOM}};
  field_stack_4_field_type_27_sub_class_id = _RAND_483[15:0];
  _RAND_484 = {1{`RANDOM}};
  field_stack_4_field_type_28_is_repeated = _RAND_484[0:0];
  _RAND_485 = {1{`RANDOM}};
  field_stack_4_field_type_28_field_type = _RAND_485[4:0];
  _RAND_486 = {1{`RANDOM}};
  field_stack_4_field_type_28_sub_class_id = _RAND_486[15:0];
  _RAND_487 = {1{`RANDOM}};
  field_stack_4_field_type_29_is_repeated = _RAND_487[0:0];
  _RAND_488 = {1{`RANDOM}};
  field_stack_4_field_type_29_field_type = _RAND_488[4:0];
  _RAND_489 = {1{`RANDOM}};
  field_stack_4_field_type_29_sub_class_id = _RAND_489[15:0];
  _RAND_490 = {1{`RANDOM}};
  field_stack_4_field_type_30_is_repeated = _RAND_490[0:0];
  _RAND_491 = {1{`RANDOM}};
  field_stack_4_field_type_30_field_type = _RAND_491[4:0];
  _RAND_492 = {1{`RANDOM}};
  field_stack_4_field_type_30_sub_class_id = _RAND_492[15:0];
  _RAND_493 = {1{`RANDOM}};
  field_stack_4_field_type_31_is_repeated = _RAND_493[0:0];
  _RAND_494 = {1{`RANDOM}};
  field_stack_4_field_type_31_field_type = _RAND_494[4:0];
  _RAND_495 = {1{`RANDOM}};
  field_stack_4_field_type_31_sub_class_id = _RAND_495[15:0];
  _RAND_496 = {1{`RANDOM}};
  field_stack_4_field_type_32_is_repeated = _RAND_496[0:0];
  _RAND_497 = {1{`RANDOM}};
  field_stack_4_field_type_32_field_type = _RAND_497[4:0];
  _RAND_498 = {1{`RANDOM}};
  field_stack_4_field_type_32_sub_class_id = _RAND_498[15:0];
  _RAND_499 = {1{`RANDOM}};
  field_stack_5_field_type_0_is_repeated = _RAND_499[0:0];
  _RAND_500 = {1{`RANDOM}};
  field_stack_5_field_type_0_field_type = _RAND_500[4:0];
  _RAND_501 = {1{`RANDOM}};
  field_stack_5_field_type_0_sub_class_id = _RAND_501[15:0];
  _RAND_502 = {1{`RANDOM}};
  field_stack_5_field_type_1_is_repeated = _RAND_502[0:0];
  _RAND_503 = {1{`RANDOM}};
  field_stack_5_field_type_1_field_type = _RAND_503[4:0];
  _RAND_504 = {1{`RANDOM}};
  field_stack_5_field_type_1_sub_class_id = _RAND_504[15:0];
  _RAND_505 = {1{`RANDOM}};
  field_stack_5_field_type_2_is_repeated = _RAND_505[0:0];
  _RAND_506 = {1{`RANDOM}};
  field_stack_5_field_type_2_field_type = _RAND_506[4:0];
  _RAND_507 = {1{`RANDOM}};
  field_stack_5_field_type_2_sub_class_id = _RAND_507[15:0];
  _RAND_508 = {1{`RANDOM}};
  field_stack_5_field_type_3_is_repeated = _RAND_508[0:0];
  _RAND_509 = {1{`RANDOM}};
  field_stack_5_field_type_3_field_type = _RAND_509[4:0];
  _RAND_510 = {1{`RANDOM}};
  field_stack_5_field_type_3_sub_class_id = _RAND_510[15:0];
  _RAND_511 = {1{`RANDOM}};
  field_stack_5_field_type_4_is_repeated = _RAND_511[0:0];
  _RAND_512 = {1{`RANDOM}};
  field_stack_5_field_type_4_field_type = _RAND_512[4:0];
  _RAND_513 = {1{`RANDOM}};
  field_stack_5_field_type_4_sub_class_id = _RAND_513[15:0];
  _RAND_514 = {1{`RANDOM}};
  field_stack_5_field_type_5_is_repeated = _RAND_514[0:0];
  _RAND_515 = {1{`RANDOM}};
  field_stack_5_field_type_5_field_type = _RAND_515[4:0];
  _RAND_516 = {1{`RANDOM}};
  field_stack_5_field_type_5_sub_class_id = _RAND_516[15:0];
  _RAND_517 = {1{`RANDOM}};
  field_stack_5_field_type_6_is_repeated = _RAND_517[0:0];
  _RAND_518 = {1{`RANDOM}};
  field_stack_5_field_type_6_field_type = _RAND_518[4:0];
  _RAND_519 = {1{`RANDOM}};
  field_stack_5_field_type_6_sub_class_id = _RAND_519[15:0];
  _RAND_520 = {1{`RANDOM}};
  field_stack_5_field_type_7_is_repeated = _RAND_520[0:0];
  _RAND_521 = {1{`RANDOM}};
  field_stack_5_field_type_7_field_type = _RAND_521[4:0];
  _RAND_522 = {1{`RANDOM}};
  field_stack_5_field_type_7_sub_class_id = _RAND_522[15:0];
  _RAND_523 = {1{`RANDOM}};
  field_stack_5_field_type_8_is_repeated = _RAND_523[0:0];
  _RAND_524 = {1{`RANDOM}};
  field_stack_5_field_type_8_field_type = _RAND_524[4:0];
  _RAND_525 = {1{`RANDOM}};
  field_stack_5_field_type_8_sub_class_id = _RAND_525[15:0];
  _RAND_526 = {1{`RANDOM}};
  field_stack_5_field_type_9_is_repeated = _RAND_526[0:0];
  _RAND_527 = {1{`RANDOM}};
  field_stack_5_field_type_9_field_type = _RAND_527[4:0];
  _RAND_528 = {1{`RANDOM}};
  field_stack_5_field_type_9_sub_class_id = _RAND_528[15:0];
  _RAND_529 = {1{`RANDOM}};
  field_stack_5_field_type_10_is_repeated = _RAND_529[0:0];
  _RAND_530 = {1{`RANDOM}};
  field_stack_5_field_type_10_field_type = _RAND_530[4:0];
  _RAND_531 = {1{`RANDOM}};
  field_stack_5_field_type_10_sub_class_id = _RAND_531[15:0];
  _RAND_532 = {1{`RANDOM}};
  field_stack_5_field_type_11_is_repeated = _RAND_532[0:0];
  _RAND_533 = {1{`RANDOM}};
  field_stack_5_field_type_11_field_type = _RAND_533[4:0];
  _RAND_534 = {1{`RANDOM}};
  field_stack_5_field_type_11_sub_class_id = _RAND_534[15:0];
  _RAND_535 = {1{`RANDOM}};
  field_stack_5_field_type_12_is_repeated = _RAND_535[0:0];
  _RAND_536 = {1{`RANDOM}};
  field_stack_5_field_type_12_field_type = _RAND_536[4:0];
  _RAND_537 = {1{`RANDOM}};
  field_stack_5_field_type_12_sub_class_id = _RAND_537[15:0];
  _RAND_538 = {1{`RANDOM}};
  field_stack_5_field_type_13_is_repeated = _RAND_538[0:0];
  _RAND_539 = {1{`RANDOM}};
  field_stack_5_field_type_13_field_type = _RAND_539[4:0];
  _RAND_540 = {1{`RANDOM}};
  field_stack_5_field_type_13_sub_class_id = _RAND_540[15:0];
  _RAND_541 = {1{`RANDOM}};
  field_stack_5_field_type_14_is_repeated = _RAND_541[0:0];
  _RAND_542 = {1{`RANDOM}};
  field_stack_5_field_type_14_field_type = _RAND_542[4:0];
  _RAND_543 = {1{`RANDOM}};
  field_stack_5_field_type_14_sub_class_id = _RAND_543[15:0];
  _RAND_544 = {1{`RANDOM}};
  field_stack_5_field_type_15_is_repeated = _RAND_544[0:0];
  _RAND_545 = {1{`RANDOM}};
  field_stack_5_field_type_15_field_type = _RAND_545[4:0];
  _RAND_546 = {1{`RANDOM}};
  field_stack_5_field_type_15_sub_class_id = _RAND_546[15:0];
  _RAND_547 = {1{`RANDOM}};
  field_stack_5_field_type_16_is_repeated = _RAND_547[0:0];
  _RAND_548 = {1{`RANDOM}};
  field_stack_5_field_type_16_field_type = _RAND_548[4:0];
  _RAND_549 = {1{`RANDOM}};
  field_stack_5_field_type_16_sub_class_id = _RAND_549[15:0];
  _RAND_550 = {1{`RANDOM}};
  field_stack_5_field_type_17_is_repeated = _RAND_550[0:0];
  _RAND_551 = {1{`RANDOM}};
  field_stack_5_field_type_17_field_type = _RAND_551[4:0];
  _RAND_552 = {1{`RANDOM}};
  field_stack_5_field_type_17_sub_class_id = _RAND_552[15:0];
  _RAND_553 = {1{`RANDOM}};
  field_stack_5_field_type_18_is_repeated = _RAND_553[0:0];
  _RAND_554 = {1{`RANDOM}};
  field_stack_5_field_type_18_field_type = _RAND_554[4:0];
  _RAND_555 = {1{`RANDOM}};
  field_stack_5_field_type_18_sub_class_id = _RAND_555[15:0];
  _RAND_556 = {1{`RANDOM}};
  field_stack_5_field_type_19_is_repeated = _RAND_556[0:0];
  _RAND_557 = {1{`RANDOM}};
  field_stack_5_field_type_19_field_type = _RAND_557[4:0];
  _RAND_558 = {1{`RANDOM}};
  field_stack_5_field_type_19_sub_class_id = _RAND_558[15:0];
  _RAND_559 = {1{`RANDOM}};
  field_stack_5_field_type_20_is_repeated = _RAND_559[0:0];
  _RAND_560 = {1{`RANDOM}};
  field_stack_5_field_type_20_field_type = _RAND_560[4:0];
  _RAND_561 = {1{`RANDOM}};
  field_stack_5_field_type_20_sub_class_id = _RAND_561[15:0];
  _RAND_562 = {1{`RANDOM}};
  field_stack_5_field_type_21_is_repeated = _RAND_562[0:0];
  _RAND_563 = {1{`RANDOM}};
  field_stack_5_field_type_21_field_type = _RAND_563[4:0];
  _RAND_564 = {1{`RANDOM}};
  field_stack_5_field_type_21_sub_class_id = _RAND_564[15:0];
  _RAND_565 = {1{`RANDOM}};
  field_stack_5_field_type_22_is_repeated = _RAND_565[0:0];
  _RAND_566 = {1{`RANDOM}};
  field_stack_5_field_type_22_field_type = _RAND_566[4:0];
  _RAND_567 = {1{`RANDOM}};
  field_stack_5_field_type_22_sub_class_id = _RAND_567[15:0];
  _RAND_568 = {1{`RANDOM}};
  field_stack_5_field_type_23_is_repeated = _RAND_568[0:0];
  _RAND_569 = {1{`RANDOM}};
  field_stack_5_field_type_23_field_type = _RAND_569[4:0];
  _RAND_570 = {1{`RANDOM}};
  field_stack_5_field_type_23_sub_class_id = _RAND_570[15:0];
  _RAND_571 = {1{`RANDOM}};
  field_stack_5_field_type_24_is_repeated = _RAND_571[0:0];
  _RAND_572 = {1{`RANDOM}};
  field_stack_5_field_type_24_field_type = _RAND_572[4:0];
  _RAND_573 = {1{`RANDOM}};
  field_stack_5_field_type_24_sub_class_id = _RAND_573[15:0];
  _RAND_574 = {1{`RANDOM}};
  field_stack_5_field_type_25_is_repeated = _RAND_574[0:0];
  _RAND_575 = {1{`RANDOM}};
  field_stack_5_field_type_25_field_type = _RAND_575[4:0];
  _RAND_576 = {1{`RANDOM}};
  field_stack_5_field_type_25_sub_class_id = _RAND_576[15:0];
  _RAND_577 = {1{`RANDOM}};
  field_stack_5_field_type_26_is_repeated = _RAND_577[0:0];
  _RAND_578 = {1{`RANDOM}};
  field_stack_5_field_type_26_field_type = _RAND_578[4:0];
  _RAND_579 = {1{`RANDOM}};
  field_stack_5_field_type_26_sub_class_id = _RAND_579[15:0];
  _RAND_580 = {1{`RANDOM}};
  field_stack_5_field_type_27_is_repeated = _RAND_580[0:0];
  _RAND_581 = {1{`RANDOM}};
  field_stack_5_field_type_27_field_type = _RAND_581[4:0];
  _RAND_582 = {1{`RANDOM}};
  field_stack_5_field_type_27_sub_class_id = _RAND_582[15:0];
  _RAND_583 = {1{`RANDOM}};
  field_stack_5_field_type_28_is_repeated = _RAND_583[0:0];
  _RAND_584 = {1{`RANDOM}};
  field_stack_5_field_type_28_field_type = _RAND_584[4:0];
  _RAND_585 = {1{`RANDOM}};
  field_stack_5_field_type_28_sub_class_id = _RAND_585[15:0];
  _RAND_586 = {1{`RANDOM}};
  field_stack_5_field_type_29_is_repeated = _RAND_586[0:0];
  _RAND_587 = {1{`RANDOM}};
  field_stack_5_field_type_29_field_type = _RAND_587[4:0];
  _RAND_588 = {1{`RANDOM}};
  field_stack_5_field_type_29_sub_class_id = _RAND_588[15:0];
  _RAND_589 = {1{`RANDOM}};
  field_stack_5_field_type_30_is_repeated = _RAND_589[0:0];
  _RAND_590 = {1{`RANDOM}};
  field_stack_5_field_type_30_field_type = _RAND_590[4:0];
  _RAND_591 = {1{`RANDOM}};
  field_stack_5_field_type_30_sub_class_id = _RAND_591[15:0];
  _RAND_592 = {1{`RANDOM}};
  field_stack_5_field_type_31_is_repeated = _RAND_592[0:0];
  _RAND_593 = {1{`RANDOM}};
  field_stack_5_field_type_31_field_type = _RAND_593[4:0];
  _RAND_594 = {1{`RANDOM}};
  field_stack_5_field_type_31_sub_class_id = _RAND_594[15:0];
  _RAND_595 = {1{`RANDOM}};
  field_stack_5_field_type_32_is_repeated = _RAND_595[0:0];
  _RAND_596 = {1{`RANDOM}};
  field_stack_5_field_type_32_field_type = _RAND_596[4:0];
  _RAND_597 = {1{`RANDOM}};
  field_stack_5_field_type_32_sub_class_id = _RAND_597[15:0];
  _RAND_598 = {1{`RANDOM}};
  field_stack_6_field_type_0_is_repeated = _RAND_598[0:0];
  _RAND_599 = {1{`RANDOM}};
  field_stack_6_field_type_0_field_type = _RAND_599[4:0];
  _RAND_600 = {1{`RANDOM}};
  field_stack_6_field_type_0_sub_class_id = _RAND_600[15:0];
  _RAND_601 = {1{`RANDOM}};
  field_stack_6_field_type_1_is_repeated = _RAND_601[0:0];
  _RAND_602 = {1{`RANDOM}};
  field_stack_6_field_type_1_field_type = _RAND_602[4:0];
  _RAND_603 = {1{`RANDOM}};
  field_stack_6_field_type_1_sub_class_id = _RAND_603[15:0];
  _RAND_604 = {1{`RANDOM}};
  field_stack_6_field_type_2_is_repeated = _RAND_604[0:0];
  _RAND_605 = {1{`RANDOM}};
  field_stack_6_field_type_2_field_type = _RAND_605[4:0];
  _RAND_606 = {1{`RANDOM}};
  field_stack_6_field_type_2_sub_class_id = _RAND_606[15:0];
  _RAND_607 = {1{`RANDOM}};
  field_stack_6_field_type_3_is_repeated = _RAND_607[0:0];
  _RAND_608 = {1{`RANDOM}};
  field_stack_6_field_type_3_field_type = _RAND_608[4:0];
  _RAND_609 = {1{`RANDOM}};
  field_stack_6_field_type_3_sub_class_id = _RAND_609[15:0];
  _RAND_610 = {1{`RANDOM}};
  field_stack_6_field_type_4_is_repeated = _RAND_610[0:0];
  _RAND_611 = {1{`RANDOM}};
  field_stack_6_field_type_4_field_type = _RAND_611[4:0];
  _RAND_612 = {1{`RANDOM}};
  field_stack_6_field_type_4_sub_class_id = _RAND_612[15:0];
  _RAND_613 = {1{`RANDOM}};
  field_stack_6_field_type_5_is_repeated = _RAND_613[0:0];
  _RAND_614 = {1{`RANDOM}};
  field_stack_6_field_type_5_field_type = _RAND_614[4:0];
  _RAND_615 = {1{`RANDOM}};
  field_stack_6_field_type_5_sub_class_id = _RAND_615[15:0];
  _RAND_616 = {1{`RANDOM}};
  field_stack_6_field_type_6_is_repeated = _RAND_616[0:0];
  _RAND_617 = {1{`RANDOM}};
  field_stack_6_field_type_6_field_type = _RAND_617[4:0];
  _RAND_618 = {1{`RANDOM}};
  field_stack_6_field_type_6_sub_class_id = _RAND_618[15:0];
  _RAND_619 = {1{`RANDOM}};
  field_stack_6_field_type_7_is_repeated = _RAND_619[0:0];
  _RAND_620 = {1{`RANDOM}};
  field_stack_6_field_type_7_field_type = _RAND_620[4:0];
  _RAND_621 = {1{`RANDOM}};
  field_stack_6_field_type_7_sub_class_id = _RAND_621[15:0];
  _RAND_622 = {1{`RANDOM}};
  field_stack_6_field_type_8_is_repeated = _RAND_622[0:0];
  _RAND_623 = {1{`RANDOM}};
  field_stack_6_field_type_8_field_type = _RAND_623[4:0];
  _RAND_624 = {1{`RANDOM}};
  field_stack_6_field_type_8_sub_class_id = _RAND_624[15:0];
  _RAND_625 = {1{`RANDOM}};
  field_stack_6_field_type_9_is_repeated = _RAND_625[0:0];
  _RAND_626 = {1{`RANDOM}};
  field_stack_6_field_type_9_field_type = _RAND_626[4:0];
  _RAND_627 = {1{`RANDOM}};
  field_stack_6_field_type_9_sub_class_id = _RAND_627[15:0];
  _RAND_628 = {1{`RANDOM}};
  field_stack_6_field_type_10_is_repeated = _RAND_628[0:0];
  _RAND_629 = {1{`RANDOM}};
  field_stack_6_field_type_10_field_type = _RAND_629[4:0];
  _RAND_630 = {1{`RANDOM}};
  field_stack_6_field_type_10_sub_class_id = _RAND_630[15:0];
  _RAND_631 = {1{`RANDOM}};
  field_stack_6_field_type_11_is_repeated = _RAND_631[0:0];
  _RAND_632 = {1{`RANDOM}};
  field_stack_6_field_type_11_field_type = _RAND_632[4:0];
  _RAND_633 = {1{`RANDOM}};
  field_stack_6_field_type_11_sub_class_id = _RAND_633[15:0];
  _RAND_634 = {1{`RANDOM}};
  field_stack_6_field_type_12_is_repeated = _RAND_634[0:0];
  _RAND_635 = {1{`RANDOM}};
  field_stack_6_field_type_12_field_type = _RAND_635[4:0];
  _RAND_636 = {1{`RANDOM}};
  field_stack_6_field_type_12_sub_class_id = _RAND_636[15:0];
  _RAND_637 = {1{`RANDOM}};
  field_stack_6_field_type_13_is_repeated = _RAND_637[0:0];
  _RAND_638 = {1{`RANDOM}};
  field_stack_6_field_type_13_field_type = _RAND_638[4:0];
  _RAND_639 = {1{`RANDOM}};
  field_stack_6_field_type_13_sub_class_id = _RAND_639[15:0];
  _RAND_640 = {1{`RANDOM}};
  field_stack_6_field_type_14_is_repeated = _RAND_640[0:0];
  _RAND_641 = {1{`RANDOM}};
  field_stack_6_field_type_14_field_type = _RAND_641[4:0];
  _RAND_642 = {1{`RANDOM}};
  field_stack_6_field_type_14_sub_class_id = _RAND_642[15:0];
  _RAND_643 = {1{`RANDOM}};
  field_stack_6_field_type_15_is_repeated = _RAND_643[0:0];
  _RAND_644 = {1{`RANDOM}};
  field_stack_6_field_type_15_field_type = _RAND_644[4:0];
  _RAND_645 = {1{`RANDOM}};
  field_stack_6_field_type_15_sub_class_id = _RAND_645[15:0];
  _RAND_646 = {1{`RANDOM}};
  field_stack_6_field_type_16_is_repeated = _RAND_646[0:0];
  _RAND_647 = {1{`RANDOM}};
  field_stack_6_field_type_16_field_type = _RAND_647[4:0];
  _RAND_648 = {1{`RANDOM}};
  field_stack_6_field_type_16_sub_class_id = _RAND_648[15:0];
  _RAND_649 = {1{`RANDOM}};
  field_stack_6_field_type_17_is_repeated = _RAND_649[0:0];
  _RAND_650 = {1{`RANDOM}};
  field_stack_6_field_type_17_field_type = _RAND_650[4:0];
  _RAND_651 = {1{`RANDOM}};
  field_stack_6_field_type_17_sub_class_id = _RAND_651[15:0];
  _RAND_652 = {1{`RANDOM}};
  field_stack_6_field_type_18_is_repeated = _RAND_652[0:0];
  _RAND_653 = {1{`RANDOM}};
  field_stack_6_field_type_18_field_type = _RAND_653[4:0];
  _RAND_654 = {1{`RANDOM}};
  field_stack_6_field_type_18_sub_class_id = _RAND_654[15:0];
  _RAND_655 = {1{`RANDOM}};
  field_stack_6_field_type_19_is_repeated = _RAND_655[0:0];
  _RAND_656 = {1{`RANDOM}};
  field_stack_6_field_type_19_field_type = _RAND_656[4:0];
  _RAND_657 = {1{`RANDOM}};
  field_stack_6_field_type_19_sub_class_id = _RAND_657[15:0];
  _RAND_658 = {1{`RANDOM}};
  field_stack_6_field_type_20_is_repeated = _RAND_658[0:0];
  _RAND_659 = {1{`RANDOM}};
  field_stack_6_field_type_20_field_type = _RAND_659[4:0];
  _RAND_660 = {1{`RANDOM}};
  field_stack_6_field_type_20_sub_class_id = _RAND_660[15:0];
  _RAND_661 = {1{`RANDOM}};
  field_stack_6_field_type_21_is_repeated = _RAND_661[0:0];
  _RAND_662 = {1{`RANDOM}};
  field_stack_6_field_type_21_field_type = _RAND_662[4:0];
  _RAND_663 = {1{`RANDOM}};
  field_stack_6_field_type_21_sub_class_id = _RAND_663[15:0];
  _RAND_664 = {1{`RANDOM}};
  field_stack_6_field_type_22_is_repeated = _RAND_664[0:0];
  _RAND_665 = {1{`RANDOM}};
  field_stack_6_field_type_22_field_type = _RAND_665[4:0];
  _RAND_666 = {1{`RANDOM}};
  field_stack_6_field_type_22_sub_class_id = _RAND_666[15:0];
  _RAND_667 = {1{`RANDOM}};
  field_stack_6_field_type_23_is_repeated = _RAND_667[0:0];
  _RAND_668 = {1{`RANDOM}};
  field_stack_6_field_type_23_field_type = _RAND_668[4:0];
  _RAND_669 = {1{`RANDOM}};
  field_stack_6_field_type_23_sub_class_id = _RAND_669[15:0];
  _RAND_670 = {1{`RANDOM}};
  field_stack_6_field_type_24_is_repeated = _RAND_670[0:0];
  _RAND_671 = {1{`RANDOM}};
  field_stack_6_field_type_24_field_type = _RAND_671[4:0];
  _RAND_672 = {1{`RANDOM}};
  field_stack_6_field_type_24_sub_class_id = _RAND_672[15:0];
  _RAND_673 = {1{`RANDOM}};
  field_stack_6_field_type_25_is_repeated = _RAND_673[0:0];
  _RAND_674 = {1{`RANDOM}};
  field_stack_6_field_type_25_field_type = _RAND_674[4:0];
  _RAND_675 = {1{`RANDOM}};
  field_stack_6_field_type_25_sub_class_id = _RAND_675[15:0];
  _RAND_676 = {1{`RANDOM}};
  field_stack_6_field_type_26_is_repeated = _RAND_676[0:0];
  _RAND_677 = {1{`RANDOM}};
  field_stack_6_field_type_26_field_type = _RAND_677[4:0];
  _RAND_678 = {1{`RANDOM}};
  field_stack_6_field_type_26_sub_class_id = _RAND_678[15:0];
  _RAND_679 = {1{`RANDOM}};
  field_stack_6_field_type_27_is_repeated = _RAND_679[0:0];
  _RAND_680 = {1{`RANDOM}};
  field_stack_6_field_type_27_field_type = _RAND_680[4:0];
  _RAND_681 = {1{`RANDOM}};
  field_stack_6_field_type_27_sub_class_id = _RAND_681[15:0];
  _RAND_682 = {1{`RANDOM}};
  field_stack_6_field_type_28_is_repeated = _RAND_682[0:0];
  _RAND_683 = {1{`RANDOM}};
  field_stack_6_field_type_28_field_type = _RAND_683[4:0];
  _RAND_684 = {1{`RANDOM}};
  field_stack_6_field_type_28_sub_class_id = _RAND_684[15:0];
  _RAND_685 = {1{`RANDOM}};
  field_stack_6_field_type_29_is_repeated = _RAND_685[0:0];
  _RAND_686 = {1{`RANDOM}};
  field_stack_6_field_type_29_field_type = _RAND_686[4:0];
  _RAND_687 = {1{`RANDOM}};
  field_stack_6_field_type_29_sub_class_id = _RAND_687[15:0];
  _RAND_688 = {1{`RANDOM}};
  field_stack_6_field_type_30_is_repeated = _RAND_688[0:0];
  _RAND_689 = {1{`RANDOM}};
  field_stack_6_field_type_30_field_type = _RAND_689[4:0];
  _RAND_690 = {1{`RANDOM}};
  field_stack_6_field_type_30_sub_class_id = _RAND_690[15:0];
  _RAND_691 = {1{`RANDOM}};
  field_stack_6_field_type_31_is_repeated = _RAND_691[0:0];
  _RAND_692 = {1{`RANDOM}};
  field_stack_6_field_type_31_field_type = _RAND_692[4:0];
  _RAND_693 = {1{`RANDOM}};
  field_stack_6_field_type_31_sub_class_id = _RAND_693[15:0];
  _RAND_694 = {1{`RANDOM}};
  field_stack_6_field_type_32_is_repeated = _RAND_694[0:0];
  _RAND_695 = {1{`RANDOM}};
  field_stack_6_field_type_32_field_type = _RAND_695[4:0];
  _RAND_696 = {1{`RANDOM}};
  field_stack_6_field_type_32_sub_class_id = _RAND_696[15:0];
  _RAND_697 = {1{`RANDOM}};
  field_stack_7_field_type_0_is_repeated = _RAND_697[0:0];
  _RAND_698 = {1{`RANDOM}};
  field_stack_7_field_type_0_field_type = _RAND_698[4:0];
  _RAND_699 = {1{`RANDOM}};
  field_stack_7_field_type_0_sub_class_id = _RAND_699[15:0];
  _RAND_700 = {1{`RANDOM}};
  field_stack_7_field_type_1_is_repeated = _RAND_700[0:0];
  _RAND_701 = {1{`RANDOM}};
  field_stack_7_field_type_1_field_type = _RAND_701[4:0];
  _RAND_702 = {1{`RANDOM}};
  field_stack_7_field_type_1_sub_class_id = _RAND_702[15:0];
  _RAND_703 = {1{`RANDOM}};
  field_stack_7_field_type_2_is_repeated = _RAND_703[0:0];
  _RAND_704 = {1{`RANDOM}};
  field_stack_7_field_type_2_field_type = _RAND_704[4:0];
  _RAND_705 = {1{`RANDOM}};
  field_stack_7_field_type_2_sub_class_id = _RAND_705[15:0];
  _RAND_706 = {1{`RANDOM}};
  field_stack_7_field_type_3_is_repeated = _RAND_706[0:0];
  _RAND_707 = {1{`RANDOM}};
  field_stack_7_field_type_3_field_type = _RAND_707[4:0];
  _RAND_708 = {1{`RANDOM}};
  field_stack_7_field_type_3_sub_class_id = _RAND_708[15:0];
  _RAND_709 = {1{`RANDOM}};
  field_stack_7_field_type_4_is_repeated = _RAND_709[0:0];
  _RAND_710 = {1{`RANDOM}};
  field_stack_7_field_type_4_field_type = _RAND_710[4:0];
  _RAND_711 = {1{`RANDOM}};
  field_stack_7_field_type_4_sub_class_id = _RAND_711[15:0];
  _RAND_712 = {1{`RANDOM}};
  field_stack_7_field_type_5_is_repeated = _RAND_712[0:0];
  _RAND_713 = {1{`RANDOM}};
  field_stack_7_field_type_5_field_type = _RAND_713[4:0];
  _RAND_714 = {1{`RANDOM}};
  field_stack_7_field_type_5_sub_class_id = _RAND_714[15:0];
  _RAND_715 = {1{`RANDOM}};
  field_stack_7_field_type_6_is_repeated = _RAND_715[0:0];
  _RAND_716 = {1{`RANDOM}};
  field_stack_7_field_type_6_field_type = _RAND_716[4:0];
  _RAND_717 = {1{`RANDOM}};
  field_stack_7_field_type_6_sub_class_id = _RAND_717[15:0];
  _RAND_718 = {1{`RANDOM}};
  field_stack_7_field_type_7_is_repeated = _RAND_718[0:0];
  _RAND_719 = {1{`RANDOM}};
  field_stack_7_field_type_7_field_type = _RAND_719[4:0];
  _RAND_720 = {1{`RANDOM}};
  field_stack_7_field_type_7_sub_class_id = _RAND_720[15:0];
  _RAND_721 = {1{`RANDOM}};
  field_stack_7_field_type_8_is_repeated = _RAND_721[0:0];
  _RAND_722 = {1{`RANDOM}};
  field_stack_7_field_type_8_field_type = _RAND_722[4:0];
  _RAND_723 = {1{`RANDOM}};
  field_stack_7_field_type_8_sub_class_id = _RAND_723[15:0];
  _RAND_724 = {1{`RANDOM}};
  field_stack_7_field_type_9_is_repeated = _RAND_724[0:0];
  _RAND_725 = {1{`RANDOM}};
  field_stack_7_field_type_9_field_type = _RAND_725[4:0];
  _RAND_726 = {1{`RANDOM}};
  field_stack_7_field_type_9_sub_class_id = _RAND_726[15:0];
  _RAND_727 = {1{`RANDOM}};
  field_stack_7_field_type_10_is_repeated = _RAND_727[0:0];
  _RAND_728 = {1{`RANDOM}};
  field_stack_7_field_type_10_field_type = _RAND_728[4:0];
  _RAND_729 = {1{`RANDOM}};
  field_stack_7_field_type_10_sub_class_id = _RAND_729[15:0];
  _RAND_730 = {1{`RANDOM}};
  field_stack_7_field_type_11_is_repeated = _RAND_730[0:0];
  _RAND_731 = {1{`RANDOM}};
  field_stack_7_field_type_11_field_type = _RAND_731[4:0];
  _RAND_732 = {1{`RANDOM}};
  field_stack_7_field_type_11_sub_class_id = _RAND_732[15:0];
  _RAND_733 = {1{`RANDOM}};
  field_stack_7_field_type_12_is_repeated = _RAND_733[0:0];
  _RAND_734 = {1{`RANDOM}};
  field_stack_7_field_type_12_field_type = _RAND_734[4:0];
  _RAND_735 = {1{`RANDOM}};
  field_stack_7_field_type_12_sub_class_id = _RAND_735[15:0];
  _RAND_736 = {1{`RANDOM}};
  field_stack_7_field_type_13_is_repeated = _RAND_736[0:0];
  _RAND_737 = {1{`RANDOM}};
  field_stack_7_field_type_13_field_type = _RAND_737[4:0];
  _RAND_738 = {1{`RANDOM}};
  field_stack_7_field_type_13_sub_class_id = _RAND_738[15:0];
  _RAND_739 = {1{`RANDOM}};
  field_stack_7_field_type_14_is_repeated = _RAND_739[0:0];
  _RAND_740 = {1{`RANDOM}};
  field_stack_7_field_type_14_field_type = _RAND_740[4:0];
  _RAND_741 = {1{`RANDOM}};
  field_stack_7_field_type_14_sub_class_id = _RAND_741[15:0];
  _RAND_742 = {1{`RANDOM}};
  field_stack_7_field_type_15_is_repeated = _RAND_742[0:0];
  _RAND_743 = {1{`RANDOM}};
  field_stack_7_field_type_15_field_type = _RAND_743[4:0];
  _RAND_744 = {1{`RANDOM}};
  field_stack_7_field_type_15_sub_class_id = _RAND_744[15:0];
  _RAND_745 = {1{`RANDOM}};
  field_stack_7_field_type_16_is_repeated = _RAND_745[0:0];
  _RAND_746 = {1{`RANDOM}};
  field_stack_7_field_type_16_field_type = _RAND_746[4:0];
  _RAND_747 = {1{`RANDOM}};
  field_stack_7_field_type_16_sub_class_id = _RAND_747[15:0];
  _RAND_748 = {1{`RANDOM}};
  field_stack_7_field_type_17_is_repeated = _RAND_748[0:0];
  _RAND_749 = {1{`RANDOM}};
  field_stack_7_field_type_17_field_type = _RAND_749[4:0];
  _RAND_750 = {1{`RANDOM}};
  field_stack_7_field_type_17_sub_class_id = _RAND_750[15:0];
  _RAND_751 = {1{`RANDOM}};
  field_stack_7_field_type_18_is_repeated = _RAND_751[0:0];
  _RAND_752 = {1{`RANDOM}};
  field_stack_7_field_type_18_field_type = _RAND_752[4:0];
  _RAND_753 = {1{`RANDOM}};
  field_stack_7_field_type_18_sub_class_id = _RAND_753[15:0];
  _RAND_754 = {1{`RANDOM}};
  field_stack_7_field_type_19_is_repeated = _RAND_754[0:0];
  _RAND_755 = {1{`RANDOM}};
  field_stack_7_field_type_19_field_type = _RAND_755[4:0];
  _RAND_756 = {1{`RANDOM}};
  field_stack_7_field_type_19_sub_class_id = _RAND_756[15:0];
  _RAND_757 = {1{`RANDOM}};
  field_stack_7_field_type_20_is_repeated = _RAND_757[0:0];
  _RAND_758 = {1{`RANDOM}};
  field_stack_7_field_type_20_field_type = _RAND_758[4:0];
  _RAND_759 = {1{`RANDOM}};
  field_stack_7_field_type_20_sub_class_id = _RAND_759[15:0];
  _RAND_760 = {1{`RANDOM}};
  field_stack_7_field_type_21_is_repeated = _RAND_760[0:0];
  _RAND_761 = {1{`RANDOM}};
  field_stack_7_field_type_21_field_type = _RAND_761[4:0];
  _RAND_762 = {1{`RANDOM}};
  field_stack_7_field_type_21_sub_class_id = _RAND_762[15:0];
  _RAND_763 = {1{`RANDOM}};
  field_stack_7_field_type_22_is_repeated = _RAND_763[0:0];
  _RAND_764 = {1{`RANDOM}};
  field_stack_7_field_type_22_field_type = _RAND_764[4:0];
  _RAND_765 = {1{`RANDOM}};
  field_stack_7_field_type_22_sub_class_id = _RAND_765[15:0];
  _RAND_766 = {1{`RANDOM}};
  field_stack_7_field_type_23_is_repeated = _RAND_766[0:0];
  _RAND_767 = {1{`RANDOM}};
  field_stack_7_field_type_23_field_type = _RAND_767[4:0];
  _RAND_768 = {1{`RANDOM}};
  field_stack_7_field_type_23_sub_class_id = _RAND_768[15:0];
  _RAND_769 = {1{`RANDOM}};
  field_stack_7_field_type_24_is_repeated = _RAND_769[0:0];
  _RAND_770 = {1{`RANDOM}};
  field_stack_7_field_type_24_field_type = _RAND_770[4:0];
  _RAND_771 = {1{`RANDOM}};
  field_stack_7_field_type_24_sub_class_id = _RAND_771[15:0];
  _RAND_772 = {1{`RANDOM}};
  field_stack_7_field_type_25_is_repeated = _RAND_772[0:0];
  _RAND_773 = {1{`RANDOM}};
  field_stack_7_field_type_25_field_type = _RAND_773[4:0];
  _RAND_774 = {1{`RANDOM}};
  field_stack_7_field_type_25_sub_class_id = _RAND_774[15:0];
  _RAND_775 = {1{`RANDOM}};
  field_stack_7_field_type_26_is_repeated = _RAND_775[0:0];
  _RAND_776 = {1{`RANDOM}};
  field_stack_7_field_type_26_field_type = _RAND_776[4:0];
  _RAND_777 = {1{`RANDOM}};
  field_stack_7_field_type_26_sub_class_id = _RAND_777[15:0];
  _RAND_778 = {1{`RANDOM}};
  field_stack_7_field_type_27_is_repeated = _RAND_778[0:0];
  _RAND_779 = {1{`RANDOM}};
  field_stack_7_field_type_27_field_type = _RAND_779[4:0];
  _RAND_780 = {1{`RANDOM}};
  field_stack_7_field_type_27_sub_class_id = _RAND_780[15:0];
  _RAND_781 = {1{`RANDOM}};
  field_stack_7_field_type_28_is_repeated = _RAND_781[0:0];
  _RAND_782 = {1{`RANDOM}};
  field_stack_7_field_type_28_field_type = _RAND_782[4:0];
  _RAND_783 = {1{`RANDOM}};
  field_stack_7_field_type_28_sub_class_id = _RAND_783[15:0];
  _RAND_784 = {1{`RANDOM}};
  field_stack_7_field_type_29_is_repeated = _RAND_784[0:0];
  _RAND_785 = {1{`RANDOM}};
  field_stack_7_field_type_29_field_type = _RAND_785[4:0];
  _RAND_786 = {1{`RANDOM}};
  field_stack_7_field_type_29_sub_class_id = _RAND_786[15:0];
  _RAND_787 = {1{`RANDOM}};
  field_stack_7_field_type_30_is_repeated = _RAND_787[0:0];
  _RAND_788 = {1{`RANDOM}};
  field_stack_7_field_type_30_field_type = _RAND_788[4:0];
  _RAND_789 = {1{`RANDOM}};
  field_stack_7_field_type_30_sub_class_id = _RAND_789[15:0];
  _RAND_790 = {1{`RANDOM}};
  field_stack_7_field_type_31_is_repeated = _RAND_790[0:0];
  _RAND_791 = {1{`RANDOM}};
  field_stack_7_field_type_31_field_type = _RAND_791[4:0];
  _RAND_792 = {1{`RANDOM}};
  field_stack_7_field_type_31_sub_class_id = _RAND_792[15:0];
  _RAND_793 = {1{`RANDOM}};
  field_stack_7_field_type_32_is_repeated = _RAND_793[0:0];
  _RAND_794 = {1{`RANDOM}};
  field_stack_7_field_type_32_field_type = _RAND_794[4:0];
  _RAND_795 = {1{`RANDOM}};
  field_stack_7_field_type_32_sub_class_id = _RAND_795[15:0];
  _RAND_796 = {1{`RANDOM}};
  field_stack_8_field_type_0_is_repeated = _RAND_796[0:0];
  _RAND_797 = {1{`RANDOM}};
  field_stack_8_field_type_0_field_type = _RAND_797[4:0];
  _RAND_798 = {1{`RANDOM}};
  field_stack_8_field_type_0_sub_class_id = _RAND_798[15:0];
  _RAND_799 = {1{`RANDOM}};
  field_stack_8_field_type_1_is_repeated = _RAND_799[0:0];
  _RAND_800 = {1{`RANDOM}};
  field_stack_8_field_type_1_field_type = _RAND_800[4:0];
  _RAND_801 = {1{`RANDOM}};
  field_stack_8_field_type_1_sub_class_id = _RAND_801[15:0];
  _RAND_802 = {1{`RANDOM}};
  field_stack_8_field_type_2_is_repeated = _RAND_802[0:0];
  _RAND_803 = {1{`RANDOM}};
  field_stack_8_field_type_2_field_type = _RAND_803[4:0];
  _RAND_804 = {1{`RANDOM}};
  field_stack_8_field_type_2_sub_class_id = _RAND_804[15:0];
  _RAND_805 = {1{`RANDOM}};
  field_stack_8_field_type_3_is_repeated = _RAND_805[0:0];
  _RAND_806 = {1{`RANDOM}};
  field_stack_8_field_type_3_field_type = _RAND_806[4:0];
  _RAND_807 = {1{`RANDOM}};
  field_stack_8_field_type_3_sub_class_id = _RAND_807[15:0];
  _RAND_808 = {1{`RANDOM}};
  field_stack_8_field_type_4_is_repeated = _RAND_808[0:0];
  _RAND_809 = {1{`RANDOM}};
  field_stack_8_field_type_4_field_type = _RAND_809[4:0];
  _RAND_810 = {1{`RANDOM}};
  field_stack_8_field_type_4_sub_class_id = _RAND_810[15:0];
  _RAND_811 = {1{`RANDOM}};
  field_stack_8_field_type_5_is_repeated = _RAND_811[0:0];
  _RAND_812 = {1{`RANDOM}};
  field_stack_8_field_type_5_field_type = _RAND_812[4:0];
  _RAND_813 = {1{`RANDOM}};
  field_stack_8_field_type_5_sub_class_id = _RAND_813[15:0];
  _RAND_814 = {1{`RANDOM}};
  field_stack_8_field_type_6_is_repeated = _RAND_814[0:0];
  _RAND_815 = {1{`RANDOM}};
  field_stack_8_field_type_6_field_type = _RAND_815[4:0];
  _RAND_816 = {1{`RANDOM}};
  field_stack_8_field_type_6_sub_class_id = _RAND_816[15:0];
  _RAND_817 = {1{`RANDOM}};
  field_stack_8_field_type_7_is_repeated = _RAND_817[0:0];
  _RAND_818 = {1{`RANDOM}};
  field_stack_8_field_type_7_field_type = _RAND_818[4:0];
  _RAND_819 = {1{`RANDOM}};
  field_stack_8_field_type_7_sub_class_id = _RAND_819[15:0];
  _RAND_820 = {1{`RANDOM}};
  field_stack_8_field_type_8_is_repeated = _RAND_820[0:0];
  _RAND_821 = {1{`RANDOM}};
  field_stack_8_field_type_8_field_type = _RAND_821[4:0];
  _RAND_822 = {1{`RANDOM}};
  field_stack_8_field_type_8_sub_class_id = _RAND_822[15:0];
  _RAND_823 = {1{`RANDOM}};
  field_stack_8_field_type_9_is_repeated = _RAND_823[0:0];
  _RAND_824 = {1{`RANDOM}};
  field_stack_8_field_type_9_field_type = _RAND_824[4:0];
  _RAND_825 = {1{`RANDOM}};
  field_stack_8_field_type_9_sub_class_id = _RAND_825[15:0];
  _RAND_826 = {1{`RANDOM}};
  field_stack_8_field_type_10_is_repeated = _RAND_826[0:0];
  _RAND_827 = {1{`RANDOM}};
  field_stack_8_field_type_10_field_type = _RAND_827[4:0];
  _RAND_828 = {1{`RANDOM}};
  field_stack_8_field_type_10_sub_class_id = _RAND_828[15:0];
  _RAND_829 = {1{`RANDOM}};
  field_stack_8_field_type_11_is_repeated = _RAND_829[0:0];
  _RAND_830 = {1{`RANDOM}};
  field_stack_8_field_type_11_field_type = _RAND_830[4:0];
  _RAND_831 = {1{`RANDOM}};
  field_stack_8_field_type_11_sub_class_id = _RAND_831[15:0];
  _RAND_832 = {1{`RANDOM}};
  field_stack_8_field_type_12_is_repeated = _RAND_832[0:0];
  _RAND_833 = {1{`RANDOM}};
  field_stack_8_field_type_12_field_type = _RAND_833[4:0];
  _RAND_834 = {1{`RANDOM}};
  field_stack_8_field_type_12_sub_class_id = _RAND_834[15:0];
  _RAND_835 = {1{`RANDOM}};
  field_stack_8_field_type_13_is_repeated = _RAND_835[0:0];
  _RAND_836 = {1{`RANDOM}};
  field_stack_8_field_type_13_field_type = _RAND_836[4:0];
  _RAND_837 = {1{`RANDOM}};
  field_stack_8_field_type_13_sub_class_id = _RAND_837[15:0];
  _RAND_838 = {1{`RANDOM}};
  field_stack_8_field_type_14_is_repeated = _RAND_838[0:0];
  _RAND_839 = {1{`RANDOM}};
  field_stack_8_field_type_14_field_type = _RAND_839[4:0];
  _RAND_840 = {1{`RANDOM}};
  field_stack_8_field_type_14_sub_class_id = _RAND_840[15:0];
  _RAND_841 = {1{`RANDOM}};
  field_stack_8_field_type_15_is_repeated = _RAND_841[0:0];
  _RAND_842 = {1{`RANDOM}};
  field_stack_8_field_type_15_field_type = _RAND_842[4:0];
  _RAND_843 = {1{`RANDOM}};
  field_stack_8_field_type_15_sub_class_id = _RAND_843[15:0];
  _RAND_844 = {1{`RANDOM}};
  field_stack_8_field_type_16_is_repeated = _RAND_844[0:0];
  _RAND_845 = {1{`RANDOM}};
  field_stack_8_field_type_16_field_type = _RAND_845[4:0];
  _RAND_846 = {1{`RANDOM}};
  field_stack_8_field_type_16_sub_class_id = _RAND_846[15:0];
  _RAND_847 = {1{`RANDOM}};
  field_stack_8_field_type_17_is_repeated = _RAND_847[0:0];
  _RAND_848 = {1{`RANDOM}};
  field_stack_8_field_type_17_field_type = _RAND_848[4:0];
  _RAND_849 = {1{`RANDOM}};
  field_stack_8_field_type_17_sub_class_id = _RAND_849[15:0];
  _RAND_850 = {1{`RANDOM}};
  field_stack_8_field_type_18_is_repeated = _RAND_850[0:0];
  _RAND_851 = {1{`RANDOM}};
  field_stack_8_field_type_18_field_type = _RAND_851[4:0];
  _RAND_852 = {1{`RANDOM}};
  field_stack_8_field_type_18_sub_class_id = _RAND_852[15:0];
  _RAND_853 = {1{`RANDOM}};
  field_stack_8_field_type_19_is_repeated = _RAND_853[0:0];
  _RAND_854 = {1{`RANDOM}};
  field_stack_8_field_type_19_field_type = _RAND_854[4:0];
  _RAND_855 = {1{`RANDOM}};
  field_stack_8_field_type_19_sub_class_id = _RAND_855[15:0];
  _RAND_856 = {1{`RANDOM}};
  field_stack_8_field_type_20_is_repeated = _RAND_856[0:0];
  _RAND_857 = {1{`RANDOM}};
  field_stack_8_field_type_20_field_type = _RAND_857[4:0];
  _RAND_858 = {1{`RANDOM}};
  field_stack_8_field_type_20_sub_class_id = _RAND_858[15:0];
  _RAND_859 = {1{`RANDOM}};
  field_stack_8_field_type_21_is_repeated = _RAND_859[0:0];
  _RAND_860 = {1{`RANDOM}};
  field_stack_8_field_type_21_field_type = _RAND_860[4:0];
  _RAND_861 = {1{`RANDOM}};
  field_stack_8_field_type_21_sub_class_id = _RAND_861[15:0];
  _RAND_862 = {1{`RANDOM}};
  field_stack_8_field_type_22_is_repeated = _RAND_862[0:0];
  _RAND_863 = {1{`RANDOM}};
  field_stack_8_field_type_22_field_type = _RAND_863[4:0];
  _RAND_864 = {1{`RANDOM}};
  field_stack_8_field_type_22_sub_class_id = _RAND_864[15:0];
  _RAND_865 = {1{`RANDOM}};
  field_stack_8_field_type_23_is_repeated = _RAND_865[0:0];
  _RAND_866 = {1{`RANDOM}};
  field_stack_8_field_type_23_field_type = _RAND_866[4:0];
  _RAND_867 = {1{`RANDOM}};
  field_stack_8_field_type_23_sub_class_id = _RAND_867[15:0];
  _RAND_868 = {1{`RANDOM}};
  field_stack_8_field_type_24_is_repeated = _RAND_868[0:0];
  _RAND_869 = {1{`RANDOM}};
  field_stack_8_field_type_24_field_type = _RAND_869[4:0];
  _RAND_870 = {1{`RANDOM}};
  field_stack_8_field_type_24_sub_class_id = _RAND_870[15:0];
  _RAND_871 = {1{`RANDOM}};
  field_stack_8_field_type_25_is_repeated = _RAND_871[0:0];
  _RAND_872 = {1{`RANDOM}};
  field_stack_8_field_type_25_field_type = _RAND_872[4:0];
  _RAND_873 = {1{`RANDOM}};
  field_stack_8_field_type_25_sub_class_id = _RAND_873[15:0];
  _RAND_874 = {1{`RANDOM}};
  field_stack_8_field_type_26_is_repeated = _RAND_874[0:0];
  _RAND_875 = {1{`RANDOM}};
  field_stack_8_field_type_26_field_type = _RAND_875[4:0];
  _RAND_876 = {1{`RANDOM}};
  field_stack_8_field_type_26_sub_class_id = _RAND_876[15:0];
  _RAND_877 = {1{`RANDOM}};
  field_stack_8_field_type_27_is_repeated = _RAND_877[0:0];
  _RAND_878 = {1{`RANDOM}};
  field_stack_8_field_type_27_field_type = _RAND_878[4:0];
  _RAND_879 = {1{`RANDOM}};
  field_stack_8_field_type_27_sub_class_id = _RAND_879[15:0];
  _RAND_880 = {1{`RANDOM}};
  field_stack_8_field_type_28_is_repeated = _RAND_880[0:0];
  _RAND_881 = {1{`RANDOM}};
  field_stack_8_field_type_28_field_type = _RAND_881[4:0];
  _RAND_882 = {1{`RANDOM}};
  field_stack_8_field_type_28_sub_class_id = _RAND_882[15:0];
  _RAND_883 = {1{`RANDOM}};
  field_stack_8_field_type_29_is_repeated = _RAND_883[0:0];
  _RAND_884 = {1{`RANDOM}};
  field_stack_8_field_type_29_field_type = _RAND_884[4:0];
  _RAND_885 = {1{`RANDOM}};
  field_stack_8_field_type_29_sub_class_id = _RAND_885[15:0];
  _RAND_886 = {1{`RANDOM}};
  field_stack_8_field_type_30_is_repeated = _RAND_886[0:0];
  _RAND_887 = {1{`RANDOM}};
  field_stack_8_field_type_30_field_type = _RAND_887[4:0];
  _RAND_888 = {1{`RANDOM}};
  field_stack_8_field_type_30_sub_class_id = _RAND_888[15:0];
  _RAND_889 = {1{`RANDOM}};
  field_stack_8_field_type_31_is_repeated = _RAND_889[0:0];
  _RAND_890 = {1{`RANDOM}};
  field_stack_8_field_type_31_field_type = _RAND_890[4:0];
  _RAND_891 = {1{`RANDOM}};
  field_stack_8_field_type_31_sub_class_id = _RAND_891[15:0];
  _RAND_892 = {1{`RANDOM}};
  field_stack_8_field_type_32_is_repeated = _RAND_892[0:0];
  _RAND_893 = {1{`RANDOM}};
  field_stack_8_field_type_32_field_type = _RAND_893[4:0];
  _RAND_894 = {1{`RANDOM}};
  field_stack_8_field_type_32_sub_class_id = _RAND_894[15:0];
  _RAND_895 = {1{`RANDOM}};
  field_stack_9_field_type_0_is_repeated = _RAND_895[0:0];
  _RAND_896 = {1{`RANDOM}};
  field_stack_9_field_type_0_field_type = _RAND_896[4:0];
  _RAND_897 = {1{`RANDOM}};
  field_stack_9_field_type_0_sub_class_id = _RAND_897[15:0];
  _RAND_898 = {1{`RANDOM}};
  field_stack_9_field_type_1_is_repeated = _RAND_898[0:0];
  _RAND_899 = {1{`RANDOM}};
  field_stack_9_field_type_1_field_type = _RAND_899[4:0];
  _RAND_900 = {1{`RANDOM}};
  field_stack_9_field_type_1_sub_class_id = _RAND_900[15:0];
  _RAND_901 = {1{`RANDOM}};
  field_stack_9_field_type_2_is_repeated = _RAND_901[0:0];
  _RAND_902 = {1{`RANDOM}};
  field_stack_9_field_type_2_field_type = _RAND_902[4:0];
  _RAND_903 = {1{`RANDOM}};
  field_stack_9_field_type_2_sub_class_id = _RAND_903[15:0];
  _RAND_904 = {1{`RANDOM}};
  field_stack_9_field_type_3_is_repeated = _RAND_904[0:0];
  _RAND_905 = {1{`RANDOM}};
  field_stack_9_field_type_3_field_type = _RAND_905[4:0];
  _RAND_906 = {1{`RANDOM}};
  field_stack_9_field_type_3_sub_class_id = _RAND_906[15:0];
  _RAND_907 = {1{`RANDOM}};
  field_stack_9_field_type_4_is_repeated = _RAND_907[0:0];
  _RAND_908 = {1{`RANDOM}};
  field_stack_9_field_type_4_field_type = _RAND_908[4:0];
  _RAND_909 = {1{`RANDOM}};
  field_stack_9_field_type_4_sub_class_id = _RAND_909[15:0];
  _RAND_910 = {1{`RANDOM}};
  field_stack_9_field_type_5_is_repeated = _RAND_910[0:0];
  _RAND_911 = {1{`RANDOM}};
  field_stack_9_field_type_5_field_type = _RAND_911[4:0];
  _RAND_912 = {1{`RANDOM}};
  field_stack_9_field_type_5_sub_class_id = _RAND_912[15:0];
  _RAND_913 = {1{`RANDOM}};
  field_stack_9_field_type_6_is_repeated = _RAND_913[0:0];
  _RAND_914 = {1{`RANDOM}};
  field_stack_9_field_type_6_field_type = _RAND_914[4:0];
  _RAND_915 = {1{`RANDOM}};
  field_stack_9_field_type_6_sub_class_id = _RAND_915[15:0];
  _RAND_916 = {1{`RANDOM}};
  field_stack_9_field_type_7_is_repeated = _RAND_916[0:0];
  _RAND_917 = {1{`RANDOM}};
  field_stack_9_field_type_7_field_type = _RAND_917[4:0];
  _RAND_918 = {1{`RANDOM}};
  field_stack_9_field_type_7_sub_class_id = _RAND_918[15:0];
  _RAND_919 = {1{`RANDOM}};
  field_stack_9_field_type_8_is_repeated = _RAND_919[0:0];
  _RAND_920 = {1{`RANDOM}};
  field_stack_9_field_type_8_field_type = _RAND_920[4:0];
  _RAND_921 = {1{`RANDOM}};
  field_stack_9_field_type_8_sub_class_id = _RAND_921[15:0];
  _RAND_922 = {1{`RANDOM}};
  field_stack_9_field_type_9_is_repeated = _RAND_922[0:0];
  _RAND_923 = {1{`RANDOM}};
  field_stack_9_field_type_9_field_type = _RAND_923[4:0];
  _RAND_924 = {1{`RANDOM}};
  field_stack_9_field_type_9_sub_class_id = _RAND_924[15:0];
  _RAND_925 = {1{`RANDOM}};
  field_stack_9_field_type_10_is_repeated = _RAND_925[0:0];
  _RAND_926 = {1{`RANDOM}};
  field_stack_9_field_type_10_field_type = _RAND_926[4:0];
  _RAND_927 = {1{`RANDOM}};
  field_stack_9_field_type_10_sub_class_id = _RAND_927[15:0];
  _RAND_928 = {1{`RANDOM}};
  field_stack_9_field_type_11_is_repeated = _RAND_928[0:0];
  _RAND_929 = {1{`RANDOM}};
  field_stack_9_field_type_11_field_type = _RAND_929[4:0];
  _RAND_930 = {1{`RANDOM}};
  field_stack_9_field_type_11_sub_class_id = _RAND_930[15:0];
  _RAND_931 = {1{`RANDOM}};
  field_stack_9_field_type_12_is_repeated = _RAND_931[0:0];
  _RAND_932 = {1{`RANDOM}};
  field_stack_9_field_type_12_field_type = _RAND_932[4:0];
  _RAND_933 = {1{`RANDOM}};
  field_stack_9_field_type_12_sub_class_id = _RAND_933[15:0];
  _RAND_934 = {1{`RANDOM}};
  field_stack_9_field_type_13_is_repeated = _RAND_934[0:0];
  _RAND_935 = {1{`RANDOM}};
  field_stack_9_field_type_13_field_type = _RAND_935[4:0];
  _RAND_936 = {1{`RANDOM}};
  field_stack_9_field_type_13_sub_class_id = _RAND_936[15:0];
  _RAND_937 = {1{`RANDOM}};
  field_stack_9_field_type_14_is_repeated = _RAND_937[0:0];
  _RAND_938 = {1{`RANDOM}};
  field_stack_9_field_type_14_field_type = _RAND_938[4:0];
  _RAND_939 = {1{`RANDOM}};
  field_stack_9_field_type_14_sub_class_id = _RAND_939[15:0];
  _RAND_940 = {1{`RANDOM}};
  field_stack_9_field_type_15_is_repeated = _RAND_940[0:0];
  _RAND_941 = {1{`RANDOM}};
  field_stack_9_field_type_15_field_type = _RAND_941[4:0];
  _RAND_942 = {1{`RANDOM}};
  field_stack_9_field_type_15_sub_class_id = _RAND_942[15:0];
  _RAND_943 = {1{`RANDOM}};
  field_stack_9_field_type_16_is_repeated = _RAND_943[0:0];
  _RAND_944 = {1{`RANDOM}};
  field_stack_9_field_type_16_field_type = _RAND_944[4:0];
  _RAND_945 = {1{`RANDOM}};
  field_stack_9_field_type_16_sub_class_id = _RAND_945[15:0];
  _RAND_946 = {1{`RANDOM}};
  field_stack_9_field_type_17_is_repeated = _RAND_946[0:0];
  _RAND_947 = {1{`RANDOM}};
  field_stack_9_field_type_17_field_type = _RAND_947[4:0];
  _RAND_948 = {1{`RANDOM}};
  field_stack_9_field_type_17_sub_class_id = _RAND_948[15:0];
  _RAND_949 = {1{`RANDOM}};
  field_stack_9_field_type_18_is_repeated = _RAND_949[0:0];
  _RAND_950 = {1{`RANDOM}};
  field_stack_9_field_type_18_field_type = _RAND_950[4:0];
  _RAND_951 = {1{`RANDOM}};
  field_stack_9_field_type_18_sub_class_id = _RAND_951[15:0];
  _RAND_952 = {1{`RANDOM}};
  field_stack_9_field_type_19_is_repeated = _RAND_952[0:0];
  _RAND_953 = {1{`RANDOM}};
  field_stack_9_field_type_19_field_type = _RAND_953[4:0];
  _RAND_954 = {1{`RANDOM}};
  field_stack_9_field_type_19_sub_class_id = _RAND_954[15:0];
  _RAND_955 = {1{`RANDOM}};
  field_stack_9_field_type_20_is_repeated = _RAND_955[0:0];
  _RAND_956 = {1{`RANDOM}};
  field_stack_9_field_type_20_field_type = _RAND_956[4:0];
  _RAND_957 = {1{`RANDOM}};
  field_stack_9_field_type_20_sub_class_id = _RAND_957[15:0];
  _RAND_958 = {1{`RANDOM}};
  field_stack_9_field_type_21_is_repeated = _RAND_958[0:0];
  _RAND_959 = {1{`RANDOM}};
  field_stack_9_field_type_21_field_type = _RAND_959[4:0];
  _RAND_960 = {1{`RANDOM}};
  field_stack_9_field_type_21_sub_class_id = _RAND_960[15:0];
  _RAND_961 = {1{`RANDOM}};
  field_stack_9_field_type_22_is_repeated = _RAND_961[0:0];
  _RAND_962 = {1{`RANDOM}};
  field_stack_9_field_type_22_field_type = _RAND_962[4:0];
  _RAND_963 = {1{`RANDOM}};
  field_stack_9_field_type_22_sub_class_id = _RAND_963[15:0];
  _RAND_964 = {1{`RANDOM}};
  field_stack_9_field_type_23_is_repeated = _RAND_964[0:0];
  _RAND_965 = {1{`RANDOM}};
  field_stack_9_field_type_23_field_type = _RAND_965[4:0];
  _RAND_966 = {1{`RANDOM}};
  field_stack_9_field_type_23_sub_class_id = _RAND_966[15:0];
  _RAND_967 = {1{`RANDOM}};
  field_stack_9_field_type_24_is_repeated = _RAND_967[0:0];
  _RAND_968 = {1{`RANDOM}};
  field_stack_9_field_type_24_field_type = _RAND_968[4:0];
  _RAND_969 = {1{`RANDOM}};
  field_stack_9_field_type_24_sub_class_id = _RAND_969[15:0];
  _RAND_970 = {1{`RANDOM}};
  field_stack_9_field_type_25_is_repeated = _RAND_970[0:0];
  _RAND_971 = {1{`RANDOM}};
  field_stack_9_field_type_25_field_type = _RAND_971[4:0];
  _RAND_972 = {1{`RANDOM}};
  field_stack_9_field_type_25_sub_class_id = _RAND_972[15:0];
  _RAND_973 = {1{`RANDOM}};
  field_stack_9_field_type_26_is_repeated = _RAND_973[0:0];
  _RAND_974 = {1{`RANDOM}};
  field_stack_9_field_type_26_field_type = _RAND_974[4:0];
  _RAND_975 = {1{`RANDOM}};
  field_stack_9_field_type_26_sub_class_id = _RAND_975[15:0];
  _RAND_976 = {1{`RANDOM}};
  field_stack_9_field_type_27_is_repeated = _RAND_976[0:0];
  _RAND_977 = {1{`RANDOM}};
  field_stack_9_field_type_27_field_type = _RAND_977[4:0];
  _RAND_978 = {1{`RANDOM}};
  field_stack_9_field_type_27_sub_class_id = _RAND_978[15:0];
  _RAND_979 = {1{`RANDOM}};
  field_stack_9_field_type_28_is_repeated = _RAND_979[0:0];
  _RAND_980 = {1{`RANDOM}};
  field_stack_9_field_type_28_field_type = _RAND_980[4:0];
  _RAND_981 = {1{`RANDOM}};
  field_stack_9_field_type_28_sub_class_id = _RAND_981[15:0];
  _RAND_982 = {1{`RANDOM}};
  field_stack_9_field_type_29_is_repeated = _RAND_982[0:0];
  _RAND_983 = {1{`RANDOM}};
  field_stack_9_field_type_29_field_type = _RAND_983[4:0];
  _RAND_984 = {1{`RANDOM}};
  field_stack_9_field_type_29_sub_class_id = _RAND_984[15:0];
  _RAND_985 = {1{`RANDOM}};
  field_stack_9_field_type_30_is_repeated = _RAND_985[0:0];
  _RAND_986 = {1{`RANDOM}};
  field_stack_9_field_type_30_field_type = _RAND_986[4:0];
  _RAND_987 = {1{`RANDOM}};
  field_stack_9_field_type_30_sub_class_id = _RAND_987[15:0];
  _RAND_988 = {1{`RANDOM}};
  field_stack_9_field_type_31_is_repeated = _RAND_988[0:0];
  _RAND_989 = {1{`RANDOM}};
  field_stack_9_field_type_31_field_type = _RAND_989[4:0];
  _RAND_990 = {1{`RANDOM}};
  field_stack_9_field_type_31_sub_class_id = _RAND_990[15:0];
  _RAND_991 = {1{`RANDOM}};
  field_stack_9_field_type_32_is_repeated = _RAND_991[0:0];
  _RAND_992 = {1{`RANDOM}};
  field_stack_9_field_type_32_field_type = _RAND_992[4:0];
  _RAND_993 = {1{`RANDOM}};
  field_stack_9_field_type_32_sub_class_id = _RAND_993[15:0];
  _RAND_994 = {1{`RANDOM}};
  field_stack_10_field_type_0_is_repeated = _RAND_994[0:0];
  _RAND_995 = {1{`RANDOM}};
  field_stack_10_field_type_0_field_type = _RAND_995[4:0];
  _RAND_996 = {1{`RANDOM}};
  field_stack_10_field_type_0_sub_class_id = _RAND_996[15:0];
  _RAND_997 = {1{`RANDOM}};
  field_stack_10_field_type_1_is_repeated = _RAND_997[0:0];
  _RAND_998 = {1{`RANDOM}};
  field_stack_10_field_type_1_field_type = _RAND_998[4:0];
  _RAND_999 = {1{`RANDOM}};
  field_stack_10_field_type_1_sub_class_id = _RAND_999[15:0];
  _RAND_1000 = {1{`RANDOM}};
  field_stack_10_field_type_2_is_repeated = _RAND_1000[0:0];
  _RAND_1001 = {1{`RANDOM}};
  field_stack_10_field_type_2_field_type = _RAND_1001[4:0];
  _RAND_1002 = {1{`RANDOM}};
  field_stack_10_field_type_2_sub_class_id = _RAND_1002[15:0];
  _RAND_1003 = {1{`RANDOM}};
  field_stack_10_field_type_3_is_repeated = _RAND_1003[0:0];
  _RAND_1004 = {1{`RANDOM}};
  field_stack_10_field_type_3_field_type = _RAND_1004[4:0];
  _RAND_1005 = {1{`RANDOM}};
  field_stack_10_field_type_3_sub_class_id = _RAND_1005[15:0];
  _RAND_1006 = {1{`RANDOM}};
  field_stack_10_field_type_4_is_repeated = _RAND_1006[0:0];
  _RAND_1007 = {1{`RANDOM}};
  field_stack_10_field_type_4_field_type = _RAND_1007[4:0];
  _RAND_1008 = {1{`RANDOM}};
  field_stack_10_field_type_4_sub_class_id = _RAND_1008[15:0];
  _RAND_1009 = {1{`RANDOM}};
  field_stack_10_field_type_5_is_repeated = _RAND_1009[0:0];
  _RAND_1010 = {1{`RANDOM}};
  field_stack_10_field_type_5_field_type = _RAND_1010[4:0];
  _RAND_1011 = {1{`RANDOM}};
  field_stack_10_field_type_5_sub_class_id = _RAND_1011[15:0];
  _RAND_1012 = {1{`RANDOM}};
  field_stack_10_field_type_6_is_repeated = _RAND_1012[0:0];
  _RAND_1013 = {1{`RANDOM}};
  field_stack_10_field_type_6_field_type = _RAND_1013[4:0];
  _RAND_1014 = {1{`RANDOM}};
  field_stack_10_field_type_6_sub_class_id = _RAND_1014[15:0];
  _RAND_1015 = {1{`RANDOM}};
  field_stack_10_field_type_7_is_repeated = _RAND_1015[0:0];
  _RAND_1016 = {1{`RANDOM}};
  field_stack_10_field_type_7_field_type = _RAND_1016[4:0];
  _RAND_1017 = {1{`RANDOM}};
  field_stack_10_field_type_7_sub_class_id = _RAND_1017[15:0];
  _RAND_1018 = {1{`RANDOM}};
  field_stack_10_field_type_8_is_repeated = _RAND_1018[0:0];
  _RAND_1019 = {1{`RANDOM}};
  field_stack_10_field_type_8_field_type = _RAND_1019[4:0];
  _RAND_1020 = {1{`RANDOM}};
  field_stack_10_field_type_8_sub_class_id = _RAND_1020[15:0];
  _RAND_1021 = {1{`RANDOM}};
  field_stack_10_field_type_9_is_repeated = _RAND_1021[0:0];
  _RAND_1022 = {1{`RANDOM}};
  field_stack_10_field_type_9_field_type = _RAND_1022[4:0];
  _RAND_1023 = {1{`RANDOM}};
  field_stack_10_field_type_9_sub_class_id = _RAND_1023[15:0];
  _RAND_1024 = {1{`RANDOM}};
  field_stack_10_field_type_10_is_repeated = _RAND_1024[0:0];
  _RAND_1025 = {1{`RANDOM}};
  field_stack_10_field_type_10_field_type = _RAND_1025[4:0];
  _RAND_1026 = {1{`RANDOM}};
  field_stack_10_field_type_10_sub_class_id = _RAND_1026[15:0];
  _RAND_1027 = {1{`RANDOM}};
  field_stack_10_field_type_11_is_repeated = _RAND_1027[0:0];
  _RAND_1028 = {1{`RANDOM}};
  field_stack_10_field_type_11_field_type = _RAND_1028[4:0];
  _RAND_1029 = {1{`RANDOM}};
  field_stack_10_field_type_11_sub_class_id = _RAND_1029[15:0];
  _RAND_1030 = {1{`RANDOM}};
  field_stack_10_field_type_12_is_repeated = _RAND_1030[0:0];
  _RAND_1031 = {1{`RANDOM}};
  field_stack_10_field_type_12_field_type = _RAND_1031[4:0];
  _RAND_1032 = {1{`RANDOM}};
  field_stack_10_field_type_12_sub_class_id = _RAND_1032[15:0];
  _RAND_1033 = {1{`RANDOM}};
  field_stack_10_field_type_13_is_repeated = _RAND_1033[0:0];
  _RAND_1034 = {1{`RANDOM}};
  field_stack_10_field_type_13_field_type = _RAND_1034[4:0];
  _RAND_1035 = {1{`RANDOM}};
  field_stack_10_field_type_13_sub_class_id = _RAND_1035[15:0];
  _RAND_1036 = {1{`RANDOM}};
  field_stack_10_field_type_14_is_repeated = _RAND_1036[0:0];
  _RAND_1037 = {1{`RANDOM}};
  field_stack_10_field_type_14_field_type = _RAND_1037[4:0];
  _RAND_1038 = {1{`RANDOM}};
  field_stack_10_field_type_14_sub_class_id = _RAND_1038[15:0];
  _RAND_1039 = {1{`RANDOM}};
  field_stack_10_field_type_15_is_repeated = _RAND_1039[0:0];
  _RAND_1040 = {1{`RANDOM}};
  field_stack_10_field_type_15_field_type = _RAND_1040[4:0];
  _RAND_1041 = {1{`RANDOM}};
  field_stack_10_field_type_15_sub_class_id = _RAND_1041[15:0];
  _RAND_1042 = {1{`RANDOM}};
  field_stack_10_field_type_16_is_repeated = _RAND_1042[0:0];
  _RAND_1043 = {1{`RANDOM}};
  field_stack_10_field_type_16_field_type = _RAND_1043[4:0];
  _RAND_1044 = {1{`RANDOM}};
  field_stack_10_field_type_16_sub_class_id = _RAND_1044[15:0];
  _RAND_1045 = {1{`RANDOM}};
  field_stack_10_field_type_17_is_repeated = _RAND_1045[0:0];
  _RAND_1046 = {1{`RANDOM}};
  field_stack_10_field_type_17_field_type = _RAND_1046[4:0];
  _RAND_1047 = {1{`RANDOM}};
  field_stack_10_field_type_17_sub_class_id = _RAND_1047[15:0];
  _RAND_1048 = {1{`RANDOM}};
  field_stack_10_field_type_18_is_repeated = _RAND_1048[0:0];
  _RAND_1049 = {1{`RANDOM}};
  field_stack_10_field_type_18_field_type = _RAND_1049[4:0];
  _RAND_1050 = {1{`RANDOM}};
  field_stack_10_field_type_18_sub_class_id = _RAND_1050[15:0];
  _RAND_1051 = {1{`RANDOM}};
  field_stack_10_field_type_19_is_repeated = _RAND_1051[0:0];
  _RAND_1052 = {1{`RANDOM}};
  field_stack_10_field_type_19_field_type = _RAND_1052[4:0];
  _RAND_1053 = {1{`RANDOM}};
  field_stack_10_field_type_19_sub_class_id = _RAND_1053[15:0];
  _RAND_1054 = {1{`RANDOM}};
  field_stack_10_field_type_20_is_repeated = _RAND_1054[0:0];
  _RAND_1055 = {1{`RANDOM}};
  field_stack_10_field_type_20_field_type = _RAND_1055[4:0];
  _RAND_1056 = {1{`RANDOM}};
  field_stack_10_field_type_20_sub_class_id = _RAND_1056[15:0];
  _RAND_1057 = {1{`RANDOM}};
  field_stack_10_field_type_21_is_repeated = _RAND_1057[0:0];
  _RAND_1058 = {1{`RANDOM}};
  field_stack_10_field_type_21_field_type = _RAND_1058[4:0];
  _RAND_1059 = {1{`RANDOM}};
  field_stack_10_field_type_21_sub_class_id = _RAND_1059[15:0];
  _RAND_1060 = {1{`RANDOM}};
  field_stack_10_field_type_22_is_repeated = _RAND_1060[0:0];
  _RAND_1061 = {1{`RANDOM}};
  field_stack_10_field_type_22_field_type = _RAND_1061[4:0];
  _RAND_1062 = {1{`RANDOM}};
  field_stack_10_field_type_22_sub_class_id = _RAND_1062[15:0];
  _RAND_1063 = {1{`RANDOM}};
  field_stack_10_field_type_23_is_repeated = _RAND_1063[0:0];
  _RAND_1064 = {1{`RANDOM}};
  field_stack_10_field_type_23_field_type = _RAND_1064[4:0];
  _RAND_1065 = {1{`RANDOM}};
  field_stack_10_field_type_23_sub_class_id = _RAND_1065[15:0];
  _RAND_1066 = {1{`RANDOM}};
  field_stack_10_field_type_24_is_repeated = _RAND_1066[0:0];
  _RAND_1067 = {1{`RANDOM}};
  field_stack_10_field_type_24_field_type = _RAND_1067[4:0];
  _RAND_1068 = {1{`RANDOM}};
  field_stack_10_field_type_24_sub_class_id = _RAND_1068[15:0];
  _RAND_1069 = {1{`RANDOM}};
  field_stack_10_field_type_25_is_repeated = _RAND_1069[0:0];
  _RAND_1070 = {1{`RANDOM}};
  field_stack_10_field_type_25_field_type = _RAND_1070[4:0];
  _RAND_1071 = {1{`RANDOM}};
  field_stack_10_field_type_25_sub_class_id = _RAND_1071[15:0];
  _RAND_1072 = {1{`RANDOM}};
  field_stack_10_field_type_26_is_repeated = _RAND_1072[0:0];
  _RAND_1073 = {1{`RANDOM}};
  field_stack_10_field_type_26_field_type = _RAND_1073[4:0];
  _RAND_1074 = {1{`RANDOM}};
  field_stack_10_field_type_26_sub_class_id = _RAND_1074[15:0];
  _RAND_1075 = {1{`RANDOM}};
  field_stack_10_field_type_27_is_repeated = _RAND_1075[0:0];
  _RAND_1076 = {1{`RANDOM}};
  field_stack_10_field_type_27_field_type = _RAND_1076[4:0];
  _RAND_1077 = {1{`RANDOM}};
  field_stack_10_field_type_27_sub_class_id = _RAND_1077[15:0];
  _RAND_1078 = {1{`RANDOM}};
  field_stack_10_field_type_28_is_repeated = _RAND_1078[0:0];
  _RAND_1079 = {1{`RANDOM}};
  field_stack_10_field_type_28_field_type = _RAND_1079[4:0];
  _RAND_1080 = {1{`RANDOM}};
  field_stack_10_field_type_28_sub_class_id = _RAND_1080[15:0];
  _RAND_1081 = {1{`RANDOM}};
  field_stack_10_field_type_29_is_repeated = _RAND_1081[0:0];
  _RAND_1082 = {1{`RANDOM}};
  field_stack_10_field_type_29_field_type = _RAND_1082[4:0];
  _RAND_1083 = {1{`RANDOM}};
  field_stack_10_field_type_29_sub_class_id = _RAND_1083[15:0];
  _RAND_1084 = {1{`RANDOM}};
  field_stack_10_field_type_30_is_repeated = _RAND_1084[0:0];
  _RAND_1085 = {1{`RANDOM}};
  field_stack_10_field_type_30_field_type = _RAND_1085[4:0];
  _RAND_1086 = {1{`RANDOM}};
  field_stack_10_field_type_30_sub_class_id = _RAND_1086[15:0];
  _RAND_1087 = {1{`RANDOM}};
  field_stack_10_field_type_31_is_repeated = _RAND_1087[0:0];
  _RAND_1088 = {1{`RANDOM}};
  field_stack_10_field_type_31_field_type = _RAND_1088[4:0];
  _RAND_1089 = {1{`RANDOM}};
  field_stack_10_field_type_31_sub_class_id = _RAND_1089[15:0];
  _RAND_1090 = {1{`RANDOM}};
  field_stack_10_field_type_32_is_repeated = _RAND_1090[0:0];
  _RAND_1091 = {1{`RANDOM}};
  field_stack_10_field_type_32_field_type = _RAND_1091[4:0];
  _RAND_1092 = {1{`RANDOM}};
  field_stack_10_field_type_32_sub_class_id = _RAND_1092[15:0];
  _RAND_1093 = {1{`RANDOM}};
  field_stack_11_field_type_0_is_repeated = _RAND_1093[0:0];
  _RAND_1094 = {1{`RANDOM}};
  field_stack_11_field_type_0_field_type = _RAND_1094[4:0];
  _RAND_1095 = {1{`RANDOM}};
  field_stack_11_field_type_0_sub_class_id = _RAND_1095[15:0];
  _RAND_1096 = {1{`RANDOM}};
  field_stack_11_field_type_1_is_repeated = _RAND_1096[0:0];
  _RAND_1097 = {1{`RANDOM}};
  field_stack_11_field_type_1_field_type = _RAND_1097[4:0];
  _RAND_1098 = {1{`RANDOM}};
  field_stack_11_field_type_1_sub_class_id = _RAND_1098[15:0];
  _RAND_1099 = {1{`RANDOM}};
  field_stack_11_field_type_2_is_repeated = _RAND_1099[0:0];
  _RAND_1100 = {1{`RANDOM}};
  field_stack_11_field_type_2_field_type = _RAND_1100[4:0];
  _RAND_1101 = {1{`RANDOM}};
  field_stack_11_field_type_2_sub_class_id = _RAND_1101[15:0];
  _RAND_1102 = {1{`RANDOM}};
  field_stack_11_field_type_3_is_repeated = _RAND_1102[0:0];
  _RAND_1103 = {1{`RANDOM}};
  field_stack_11_field_type_3_field_type = _RAND_1103[4:0];
  _RAND_1104 = {1{`RANDOM}};
  field_stack_11_field_type_3_sub_class_id = _RAND_1104[15:0];
  _RAND_1105 = {1{`RANDOM}};
  field_stack_11_field_type_4_is_repeated = _RAND_1105[0:0];
  _RAND_1106 = {1{`RANDOM}};
  field_stack_11_field_type_4_field_type = _RAND_1106[4:0];
  _RAND_1107 = {1{`RANDOM}};
  field_stack_11_field_type_4_sub_class_id = _RAND_1107[15:0];
  _RAND_1108 = {1{`RANDOM}};
  field_stack_11_field_type_5_is_repeated = _RAND_1108[0:0];
  _RAND_1109 = {1{`RANDOM}};
  field_stack_11_field_type_5_field_type = _RAND_1109[4:0];
  _RAND_1110 = {1{`RANDOM}};
  field_stack_11_field_type_5_sub_class_id = _RAND_1110[15:0];
  _RAND_1111 = {1{`RANDOM}};
  field_stack_11_field_type_6_is_repeated = _RAND_1111[0:0];
  _RAND_1112 = {1{`RANDOM}};
  field_stack_11_field_type_6_field_type = _RAND_1112[4:0];
  _RAND_1113 = {1{`RANDOM}};
  field_stack_11_field_type_6_sub_class_id = _RAND_1113[15:0];
  _RAND_1114 = {1{`RANDOM}};
  field_stack_11_field_type_7_is_repeated = _RAND_1114[0:0];
  _RAND_1115 = {1{`RANDOM}};
  field_stack_11_field_type_7_field_type = _RAND_1115[4:0];
  _RAND_1116 = {1{`RANDOM}};
  field_stack_11_field_type_7_sub_class_id = _RAND_1116[15:0];
  _RAND_1117 = {1{`RANDOM}};
  field_stack_11_field_type_8_is_repeated = _RAND_1117[0:0];
  _RAND_1118 = {1{`RANDOM}};
  field_stack_11_field_type_8_field_type = _RAND_1118[4:0];
  _RAND_1119 = {1{`RANDOM}};
  field_stack_11_field_type_8_sub_class_id = _RAND_1119[15:0];
  _RAND_1120 = {1{`RANDOM}};
  field_stack_11_field_type_9_is_repeated = _RAND_1120[0:0];
  _RAND_1121 = {1{`RANDOM}};
  field_stack_11_field_type_9_field_type = _RAND_1121[4:0];
  _RAND_1122 = {1{`RANDOM}};
  field_stack_11_field_type_9_sub_class_id = _RAND_1122[15:0];
  _RAND_1123 = {1{`RANDOM}};
  field_stack_11_field_type_10_is_repeated = _RAND_1123[0:0];
  _RAND_1124 = {1{`RANDOM}};
  field_stack_11_field_type_10_field_type = _RAND_1124[4:0];
  _RAND_1125 = {1{`RANDOM}};
  field_stack_11_field_type_10_sub_class_id = _RAND_1125[15:0];
  _RAND_1126 = {1{`RANDOM}};
  field_stack_11_field_type_11_is_repeated = _RAND_1126[0:0];
  _RAND_1127 = {1{`RANDOM}};
  field_stack_11_field_type_11_field_type = _RAND_1127[4:0];
  _RAND_1128 = {1{`RANDOM}};
  field_stack_11_field_type_11_sub_class_id = _RAND_1128[15:0];
  _RAND_1129 = {1{`RANDOM}};
  field_stack_11_field_type_12_is_repeated = _RAND_1129[0:0];
  _RAND_1130 = {1{`RANDOM}};
  field_stack_11_field_type_12_field_type = _RAND_1130[4:0];
  _RAND_1131 = {1{`RANDOM}};
  field_stack_11_field_type_12_sub_class_id = _RAND_1131[15:0];
  _RAND_1132 = {1{`RANDOM}};
  field_stack_11_field_type_13_is_repeated = _RAND_1132[0:0];
  _RAND_1133 = {1{`RANDOM}};
  field_stack_11_field_type_13_field_type = _RAND_1133[4:0];
  _RAND_1134 = {1{`RANDOM}};
  field_stack_11_field_type_13_sub_class_id = _RAND_1134[15:0];
  _RAND_1135 = {1{`RANDOM}};
  field_stack_11_field_type_14_is_repeated = _RAND_1135[0:0];
  _RAND_1136 = {1{`RANDOM}};
  field_stack_11_field_type_14_field_type = _RAND_1136[4:0];
  _RAND_1137 = {1{`RANDOM}};
  field_stack_11_field_type_14_sub_class_id = _RAND_1137[15:0];
  _RAND_1138 = {1{`RANDOM}};
  field_stack_11_field_type_15_is_repeated = _RAND_1138[0:0];
  _RAND_1139 = {1{`RANDOM}};
  field_stack_11_field_type_15_field_type = _RAND_1139[4:0];
  _RAND_1140 = {1{`RANDOM}};
  field_stack_11_field_type_15_sub_class_id = _RAND_1140[15:0];
  _RAND_1141 = {1{`RANDOM}};
  field_stack_11_field_type_16_is_repeated = _RAND_1141[0:0];
  _RAND_1142 = {1{`RANDOM}};
  field_stack_11_field_type_16_field_type = _RAND_1142[4:0];
  _RAND_1143 = {1{`RANDOM}};
  field_stack_11_field_type_16_sub_class_id = _RAND_1143[15:0];
  _RAND_1144 = {1{`RANDOM}};
  field_stack_11_field_type_17_is_repeated = _RAND_1144[0:0];
  _RAND_1145 = {1{`RANDOM}};
  field_stack_11_field_type_17_field_type = _RAND_1145[4:0];
  _RAND_1146 = {1{`RANDOM}};
  field_stack_11_field_type_17_sub_class_id = _RAND_1146[15:0];
  _RAND_1147 = {1{`RANDOM}};
  field_stack_11_field_type_18_is_repeated = _RAND_1147[0:0];
  _RAND_1148 = {1{`RANDOM}};
  field_stack_11_field_type_18_field_type = _RAND_1148[4:0];
  _RAND_1149 = {1{`RANDOM}};
  field_stack_11_field_type_18_sub_class_id = _RAND_1149[15:0];
  _RAND_1150 = {1{`RANDOM}};
  field_stack_11_field_type_19_is_repeated = _RAND_1150[0:0];
  _RAND_1151 = {1{`RANDOM}};
  field_stack_11_field_type_19_field_type = _RAND_1151[4:0];
  _RAND_1152 = {1{`RANDOM}};
  field_stack_11_field_type_19_sub_class_id = _RAND_1152[15:0];
  _RAND_1153 = {1{`RANDOM}};
  field_stack_11_field_type_20_is_repeated = _RAND_1153[0:0];
  _RAND_1154 = {1{`RANDOM}};
  field_stack_11_field_type_20_field_type = _RAND_1154[4:0];
  _RAND_1155 = {1{`RANDOM}};
  field_stack_11_field_type_20_sub_class_id = _RAND_1155[15:0];
  _RAND_1156 = {1{`RANDOM}};
  field_stack_11_field_type_21_is_repeated = _RAND_1156[0:0];
  _RAND_1157 = {1{`RANDOM}};
  field_stack_11_field_type_21_field_type = _RAND_1157[4:0];
  _RAND_1158 = {1{`RANDOM}};
  field_stack_11_field_type_21_sub_class_id = _RAND_1158[15:0];
  _RAND_1159 = {1{`RANDOM}};
  field_stack_11_field_type_22_is_repeated = _RAND_1159[0:0];
  _RAND_1160 = {1{`RANDOM}};
  field_stack_11_field_type_22_field_type = _RAND_1160[4:0];
  _RAND_1161 = {1{`RANDOM}};
  field_stack_11_field_type_22_sub_class_id = _RAND_1161[15:0];
  _RAND_1162 = {1{`RANDOM}};
  field_stack_11_field_type_23_is_repeated = _RAND_1162[0:0];
  _RAND_1163 = {1{`RANDOM}};
  field_stack_11_field_type_23_field_type = _RAND_1163[4:0];
  _RAND_1164 = {1{`RANDOM}};
  field_stack_11_field_type_23_sub_class_id = _RAND_1164[15:0];
  _RAND_1165 = {1{`RANDOM}};
  field_stack_11_field_type_24_is_repeated = _RAND_1165[0:0];
  _RAND_1166 = {1{`RANDOM}};
  field_stack_11_field_type_24_field_type = _RAND_1166[4:0];
  _RAND_1167 = {1{`RANDOM}};
  field_stack_11_field_type_24_sub_class_id = _RAND_1167[15:0];
  _RAND_1168 = {1{`RANDOM}};
  field_stack_11_field_type_25_is_repeated = _RAND_1168[0:0];
  _RAND_1169 = {1{`RANDOM}};
  field_stack_11_field_type_25_field_type = _RAND_1169[4:0];
  _RAND_1170 = {1{`RANDOM}};
  field_stack_11_field_type_25_sub_class_id = _RAND_1170[15:0];
  _RAND_1171 = {1{`RANDOM}};
  field_stack_11_field_type_26_is_repeated = _RAND_1171[0:0];
  _RAND_1172 = {1{`RANDOM}};
  field_stack_11_field_type_26_field_type = _RAND_1172[4:0];
  _RAND_1173 = {1{`RANDOM}};
  field_stack_11_field_type_26_sub_class_id = _RAND_1173[15:0];
  _RAND_1174 = {1{`RANDOM}};
  field_stack_11_field_type_27_is_repeated = _RAND_1174[0:0];
  _RAND_1175 = {1{`RANDOM}};
  field_stack_11_field_type_27_field_type = _RAND_1175[4:0];
  _RAND_1176 = {1{`RANDOM}};
  field_stack_11_field_type_27_sub_class_id = _RAND_1176[15:0];
  _RAND_1177 = {1{`RANDOM}};
  field_stack_11_field_type_28_is_repeated = _RAND_1177[0:0];
  _RAND_1178 = {1{`RANDOM}};
  field_stack_11_field_type_28_field_type = _RAND_1178[4:0];
  _RAND_1179 = {1{`RANDOM}};
  field_stack_11_field_type_28_sub_class_id = _RAND_1179[15:0];
  _RAND_1180 = {1{`RANDOM}};
  field_stack_11_field_type_29_is_repeated = _RAND_1180[0:0];
  _RAND_1181 = {1{`RANDOM}};
  field_stack_11_field_type_29_field_type = _RAND_1181[4:0];
  _RAND_1182 = {1{`RANDOM}};
  field_stack_11_field_type_29_sub_class_id = _RAND_1182[15:0];
  _RAND_1183 = {1{`RANDOM}};
  field_stack_11_field_type_30_is_repeated = _RAND_1183[0:0];
  _RAND_1184 = {1{`RANDOM}};
  field_stack_11_field_type_30_field_type = _RAND_1184[4:0];
  _RAND_1185 = {1{`RANDOM}};
  field_stack_11_field_type_30_sub_class_id = _RAND_1185[15:0];
  _RAND_1186 = {1{`RANDOM}};
  field_stack_11_field_type_31_is_repeated = _RAND_1186[0:0];
  _RAND_1187 = {1{`RANDOM}};
  field_stack_11_field_type_31_field_type = _RAND_1187[4:0];
  _RAND_1188 = {1{`RANDOM}};
  field_stack_11_field_type_31_sub_class_id = _RAND_1188[15:0];
  _RAND_1189 = {1{`RANDOM}};
  field_stack_11_field_type_32_is_repeated = _RAND_1189[0:0];
  _RAND_1190 = {1{`RANDOM}};
  field_stack_11_field_type_32_field_type = _RAND_1190[4:0];
  _RAND_1191 = {1{`RANDOM}};
  field_stack_11_field_type_32_sub_class_id = _RAND_1191[15:0];
  _RAND_1192 = {1{`RANDOM}};
  field_stack_12_field_type_0_is_repeated = _RAND_1192[0:0];
  _RAND_1193 = {1{`RANDOM}};
  field_stack_12_field_type_0_field_type = _RAND_1193[4:0];
  _RAND_1194 = {1{`RANDOM}};
  field_stack_12_field_type_0_sub_class_id = _RAND_1194[15:0];
  _RAND_1195 = {1{`RANDOM}};
  field_stack_12_field_type_1_is_repeated = _RAND_1195[0:0];
  _RAND_1196 = {1{`RANDOM}};
  field_stack_12_field_type_1_field_type = _RAND_1196[4:0];
  _RAND_1197 = {1{`RANDOM}};
  field_stack_12_field_type_1_sub_class_id = _RAND_1197[15:0];
  _RAND_1198 = {1{`RANDOM}};
  field_stack_12_field_type_2_is_repeated = _RAND_1198[0:0];
  _RAND_1199 = {1{`RANDOM}};
  field_stack_12_field_type_2_field_type = _RAND_1199[4:0];
  _RAND_1200 = {1{`RANDOM}};
  field_stack_12_field_type_2_sub_class_id = _RAND_1200[15:0];
  _RAND_1201 = {1{`RANDOM}};
  field_stack_12_field_type_3_is_repeated = _RAND_1201[0:0];
  _RAND_1202 = {1{`RANDOM}};
  field_stack_12_field_type_3_field_type = _RAND_1202[4:0];
  _RAND_1203 = {1{`RANDOM}};
  field_stack_12_field_type_3_sub_class_id = _RAND_1203[15:0];
  _RAND_1204 = {1{`RANDOM}};
  field_stack_12_field_type_4_is_repeated = _RAND_1204[0:0];
  _RAND_1205 = {1{`RANDOM}};
  field_stack_12_field_type_4_field_type = _RAND_1205[4:0];
  _RAND_1206 = {1{`RANDOM}};
  field_stack_12_field_type_4_sub_class_id = _RAND_1206[15:0];
  _RAND_1207 = {1{`RANDOM}};
  field_stack_12_field_type_5_is_repeated = _RAND_1207[0:0];
  _RAND_1208 = {1{`RANDOM}};
  field_stack_12_field_type_5_field_type = _RAND_1208[4:0];
  _RAND_1209 = {1{`RANDOM}};
  field_stack_12_field_type_5_sub_class_id = _RAND_1209[15:0];
  _RAND_1210 = {1{`RANDOM}};
  field_stack_12_field_type_6_is_repeated = _RAND_1210[0:0];
  _RAND_1211 = {1{`RANDOM}};
  field_stack_12_field_type_6_field_type = _RAND_1211[4:0];
  _RAND_1212 = {1{`RANDOM}};
  field_stack_12_field_type_6_sub_class_id = _RAND_1212[15:0];
  _RAND_1213 = {1{`RANDOM}};
  field_stack_12_field_type_7_is_repeated = _RAND_1213[0:0];
  _RAND_1214 = {1{`RANDOM}};
  field_stack_12_field_type_7_field_type = _RAND_1214[4:0];
  _RAND_1215 = {1{`RANDOM}};
  field_stack_12_field_type_7_sub_class_id = _RAND_1215[15:0];
  _RAND_1216 = {1{`RANDOM}};
  field_stack_12_field_type_8_is_repeated = _RAND_1216[0:0];
  _RAND_1217 = {1{`RANDOM}};
  field_stack_12_field_type_8_field_type = _RAND_1217[4:0];
  _RAND_1218 = {1{`RANDOM}};
  field_stack_12_field_type_8_sub_class_id = _RAND_1218[15:0];
  _RAND_1219 = {1{`RANDOM}};
  field_stack_12_field_type_9_is_repeated = _RAND_1219[0:0];
  _RAND_1220 = {1{`RANDOM}};
  field_stack_12_field_type_9_field_type = _RAND_1220[4:0];
  _RAND_1221 = {1{`RANDOM}};
  field_stack_12_field_type_9_sub_class_id = _RAND_1221[15:0];
  _RAND_1222 = {1{`RANDOM}};
  field_stack_12_field_type_10_is_repeated = _RAND_1222[0:0];
  _RAND_1223 = {1{`RANDOM}};
  field_stack_12_field_type_10_field_type = _RAND_1223[4:0];
  _RAND_1224 = {1{`RANDOM}};
  field_stack_12_field_type_10_sub_class_id = _RAND_1224[15:0];
  _RAND_1225 = {1{`RANDOM}};
  field_stack_12_field_type_11_is_repeated = _RAND_1225[0:0];
  _RAND_1226 = {1{`RANDOM}};
  field_stack_12_field_type_11_field_type = _RAND_1226[4:0];
  _RAND_1227 = {1{`RANDOM}};
  field_stack_12_field_type_11_sub_class_id = _RAND_1227[15:0];
  _RAND_1228 = {1{`RANDOM}};
  field_stack_12_field_type_12_is_repeated = _RAND_1228[0:0];
  _RAND_1229 = {1{`RANDOM}};
  field_stack_12_field_type_12_field_type = _RAND_1229[4:0];
  _RAND_1230 = {1{`RANDOM}};
  field_stack_12_field_type_12_sub_class_id = _RAND_1230[15:0];
  _RAND_1231 = {1{`RANDOM}};
  field_stack_12_field_type_13_is_repeated = _RAND_1231[0:0];
  _RAND_1232 = {1{`RANDOM}};
  field_stack_12_field_type_13_field_type = _RAND_1232[4:0];
  _RAND_1233 = {1{`RANDOM}};
  field_stack_12_field_type_13_sub_class_id = _RAND_1233[15:0];
  _RAND_1234 = {1{`RANDOM}};
  field_stack_12_field_type_14_is_repeated = _RAND_1234[0:0];
  _RAND_1235 = {1{`RANDOM}};
  field_stack_12_field_type_14_field_type = _RAND_1235[4:0];
  _RAND_1236 = {1{`RANDOM}};
  field_stack_12_field_type_14_sub_class_id = _RAND_1236[15:0];
  _RAND_1237 = {1{`RANDOM}};
  field_stack_12_field_type_15_is_repeated = _RAND_1237[0:0];
  _RAND_1238 = {1{`RANDOM}};
  field_stack_12_field_type_15_field_type = _RAND_1238[4:0];
  _RAND_1239 = {1{`RANDOM}};
  field_stack_12_field_type_15_sub_class_id = _RAND_1239[15:0];
  _RAND_1240 = {1{`RANDOM}};
  field_stack_12_field_type_16_is_repeated = _RAND_1240[0:0];
  _RAND_1241 = {1{`RANDOM}};
  field_stack_12_field_type_16_field_type = _RAND_1241[4:0];
  _RAND_1242 = {1{`RANDOM}};
  field_stack_12_field_type_16_sub_class_id = _RAND_1242[15:0];
  _RAND_1243 = {1{`RANDOM}};
  field_stack_12_field_type_17_is_repeated = _RAND_1243[0:0];
  _RAND_1244 = {1{`RANDOM}};
  field_stack_12_field_type_17_field_type = _RAND_1244[4:0];
  _RAND_1245 = {1{`RANDOM}};
  field_stack_12_field_type_17_sub_class_id = _RAND_1245[15:0];
  _RAND_1246 = {1{`RANDOM}};
  field_stack_12_field_type_18_is_repeated = _RAND_1246[0:0];
  _RAND_1247 = {1{`RANDOM}};
  field_stack_12_field_type_18_field_type = _RAND_1247[4:0];
  _RAND_1248 = {1{`RANDOM}};
  field_stack_12_field_type_18_sub_class_id = _RAND_1248[15:0];
  _RAND_1249 = {1{`RANDOM}};
  field_stack_12_field_type_19_is_repeated = _RAND_1249[0:0];
  _RAND_1250 = {1{`RANDOM}};
  field_stack_12_field_type_19_field_type = _RAND_1250[4:0];
  _RAND_1251 = {1{`RANDOM}};
  field_stack_12_field_type_19_sub_class_id = _RAND_1251[15:0];
  _RAND_1252 = {1{`RANDOM}};
  field_stack_12_field_type_20_is_repeated = _RAND_1252[0:0];
  _RAND_1253 = {1{`RANDOM}};
  field_stack_12_field_type_20_field_type = _RAND_1253[4:0];
  _RAND_1254 = {1{`RANDOM}};
  field_stack_12_field_type_20_sub_class_id = _RAND_1254[15:0];
  _RAND_1255 = {1{`RANDOM}};
  field_stack_12_field_type_21_is_repeated = _RAND_1255[0:0];
  _RAND_1256 = {1{`RANDOM}};
  field_stack_12_field_type_21_field_type = _RAND_1256[4:0];
  _RAND_1257 = {1{`RANDOM}};
  field_stack_12_field_type_21_sub_class_id = _RAND_1257[15:0];
  _RAND_1258 = {1{`RANDOM}};
  field_stack_12_field_type_22_is_repeated = _RAND_1258[0:0];
  _RAND_1259 = {1{`RANDOM}};
  field_stack_12_field_type_22_field_type = _RAND_1259[4:0];
  _RAND_1260 = {1{`RANDOM}};
  field_stack_12_field_type_22_sub_class_id = _RAND_1260[15:0];
  _RAND_1261 = {1{`RANDOM}};
  field_stack_12_field_type_23_is_repeated = _RAND_1261[0:0];
  _RAND_1262 = {1{`RANDOM}};
  field_stack_12_field_type_23_field_type = _RAND_1262[4:0];
  _RAND_1263 = {1{`RANDOM}};
  field_stack_12_field_type_23_sub_class_id = _RAND_1263[15:0];
  _RAND_1264 = {1{`RANDOM}};
  field_stack_12_field_type_24_is_repeated = _RAND_1264[0:0];
  _RAND_1265 = {1{`RANDOM}};
  field_stack_12_field_type_24_field_type = _RAND_1265[4:0];
  _RAND_1266 = {1{`RANDOM}};
  field_stack_12_field_type_24_sub_class_id = _RAND_1266[15:0];
  _RAND_1267 = {1{`RANDOM}};
  field_stack_12_field_type_25_is_repeated = _RAND_1267[0:0];
  _RAND_1268 = {1{`RANDOM}};
  field_stack_12_field_type_25_field_type = _RAND_1268[4:0];
  _RAND_1269 = {1{`RANDOM}};
  field_stack_12_field_type_25_sub_class_id = _RAND_1269[15:0];
  _RAND_1270 = {1{`RANDOM}};
  field_stack_12_field_type_26_is_repeated = _RAND_1270[0:0];
  _RAND_1271 = {1{`RANDOM}};
  field_stack_12_field_type_26_field_type = _RAND_1271[4:0];
  _RAND_1272 = {1{`RANDOM}};
  field_stack_12_field_type_26_sub_class_id = _RAND_1272[15:0];
  _RAND_1273 = {1{`RANDOM}};
  field_stack_12_field_type_27_is_repeated = _RAND_1273[0:0];
  _RAND_1274 = {1{`RANDOM}};
  field_stack_12_field_type_27_field_type = _RAND_1274[4:0];
  _RAND_1275 = {1{`RANDOM}};
  field_stack_12_field_type_27_sub_class_id = _RAND_1275[15:0];
  _RAND_1276 = {1{`RANDOM}};
  field_stack_12_field_type_28_is_repeated = _RAND_1276[0:0];
  _RAND_1277 = {1{`RANDOM}};
  field_stack_12_field_type_28_field_type = _RAND_1277[4:0];
  _RAND_1278 = {1{`RANDOM}};
  field_stack_12_field_type_28_sub_class_id = _RAND_1278[15:0];
  _RAND_1279 = {1{`RANDOM}};
  field_stack_12_field_type_29_is_repeated = _RAND_1279[0:0];
  _RAND_1280 = {1{`RANDOM}};
  field_stack_12_field_type_29_field_type = _RAND_1280[4:0];
  _RAND_1281 = {1{`RANDOM}};
  field_stack_12_field_type_29_sub_class_id = _RAND_1281[15:0];
  _RAND_1282 = {1{`RANDOM}};
  field_stack_12_field_type_30_is_repeated = _RAND_1282[0:0];
  _RAND_1283 = {1{`RANDOM}};
  field_stack_12_field_type_30_field_type = _RAND_1283[4:0];
  _RAND_1284 = {1{`RANDOM}};
  field_stack_12_field_type_30_sub_class_id = _RAND_1284[15:0];
  _RAND_1285 = {1{`RANDOM}};
  field_stack_12_field_type_31_is_repeated = _RAND_1285[0:0];
  _RAND_1286 = {1{`RANDOM}};
  field_stack_12_field_type_31_field_type = _RAND_1286[4:0];
  _RAND_1287 = {1{`RANDOM}};
  field_stack_12_field_type_31_sub_class_id = _RAND_1287[15:0];
  _RAND_1288 = {1{`RANDOM}};
  field_stack_12_field_type_32_is_repeated = _RAND_1288[0:0];
  _RAND_1289 = {1{`RANDOM}};
  field_stack_12_field_type_32_field_type = _RAND_1289[4:0];
  _RAND_1290 = {1{`RANDOM}};
  field_stack_12_field_type_32_sub_class_id = _RAND_1290[15:0];
  _RAND_1291 = {1{`RANDOM}};
  field_stack_13_field_type_0_is_repeated = _RAND_1291[0:0];
  _RAND_1292 = {1{`RANDOM}};
  field_stack_13_field_type_0_field_type = _RAND_1292[4:0];
  _RAND_1293 = {1{`RANDOM}};
  field_stack_13_field_type_0_sub_class_id = _RAND_1293[15:0];
  _RAND_1294 = {1{`RANDOM}};
  field_stack_13_field_type_1_is_repeated = _RAND_1294[0:0];
  _RAND_1295 = {1{`RANDOM}};
  field_stack_13_field_type_1_field_type = _RAND_1295[4:0];
  _RAND_1296 = {1{`RANDOM}};
  field_stack_13_field_type_1_sub_class_id = _RAND_1296[15:0];
  _RAND_1297 = {1{`RANDOM}};
  field_stack_13_field_type_2_is_repeated = _RAND_1297[0:0];
  _RAND_1298 = {1{`RANDOM}};
  field_stack_13_field_type_2_field_type = _RAND_1298[4:0];
  _RAND_1299 = {1{`RANDOM}};
  field_stack_13_field_type_2_sub_class_id = _RAND_1299[15:0];
  _RAND_1300 = {1{`RANDOM}};
  field_stack_13_field_type_3_is_repeated = _RAND_1300[0:0];
  _RAND_1301 = {1{`RANDOM}};
  field_stack_13_field_type_3_field_type = _RAND_1301[4:0];
  _RAND_1302 = {1{`RANDOM}};
  field_stack_13_field_type_3_sub_class_id = _RAND_1302[15:0];
  _RAND_1303 = {1{`RANDOM}};
  field_stack_13_field_type_4_is_repeated = _RAND_1303[0:0];
  _RAND_1304 = {1{`RANDOM}};
  field_stack_13_field_type_4_field_type = _RAND_1304[4:0];
  _RAND_1305 = {1{`RANDOM}};
  field_stack_13_field_type_4_sub_class_id = _RAND_1305[15:0];
  _RAND_1306 = {1{`RANDOM}};
  field_stack_13_field_type_5_is_repeated = _RAND_1306[0:0];
  _RAND_1307 = {1{`RANDOM}};
  field_stack_13_field_type_5_field_type = _RAND_1307[4:0];
  _RAND_1308 = {1{`RANDOM}};
  field_stack_13_field_type_5_sub_class_id = _RAND_1308[15:0];
  _RAND_1309 = {1{`RANDOM}};
  field_stack_13_field_type_6_is_repeated = _RAND_1309[0:0];
  _RAND_1310 = {1{`RANDOM}};
  field_stack_13_field_type_6_field_type = _RAND_1310[4:0];
  _RAND_1311 = {1{`RANDOM}};
  field_stack_13_field_type_6_sub_class_id = _RAND_1311[15:0];
  _RAND_1312 = {1{`RANDOM}};
  field_stack_13_field_type_7_is_repeated = _RAND_1312[0:0];
  _RAND_1313 = {1{`RANDOM}};
  field_stack_13_field_type_7_field_type = _RAND_1313[4:0];
  _RAND_1314 = {1{`RANDOM}};
  field_stack_13_field_type_7_sub_class_id = _RAND_1314[15:0];
  _RAND_1315 = {1{`RANDOM}};
  field_stack_13_field_type_8_is_repeated = _RAND_1315[0:0];
  _RAND_1316 = {1{`RANDOM}};
  field_stack_13_field_type_8_field_type = _RAND_1316[4:0];
  _RAND_1317 = {1{`RANDOM}};
  field_stack_13_field_type_8_sub_class_id = _RAND_1317[15:0];
  _RAND_1318 = {1{`RANDOM}};
  field_stack_13_field_type_9_is_repeated = _RAND_1318[0:0];
  _RAND_1319 = {1{`RANDOM}};
  field_stack_13_field_type_9_field_type = _RAND_1319[4:0];
  _RAND_1320 = {1{`RANDOM}};
  field_stack_13_field_type_9_sub_class_id = _RAND_1320[15:0];
  _RAND_1321 = {1{`RANDOM}};
  field_stack_13_field_type_10_is_repeated = _RAND_1321[0:0];
  _RAND_1322 = {1{`RANDOM}};
  field_stack_13_field_type_10_field_type = _RAND_1322[4:0];
  _RAND_1323 = {1{`RANDOM}};
  field_stack_13_field_type_10_sub_class_id = _RAND_1323[15:0];
  _RAND_1324 = {1{`RANDOM}};
  field_stack_13_field_type_11_is_repeated = _RAND_1324[0:0];
  _RAND_1325 = {1{`RANDOM}};
  field_stack_13_field_type_11_field_type = _RAND_1325[4:0];
  _RAND_1326 = {1{`RANDOM}};
  field_stack_13_field_type_11_sub_class_id = _RAND_1326[15:0];
  _RAND_1327 = {1{`RANDOM}};
  field_stack_13_field_type_12_is_repeated = _RAND_1327[0:0];
  _RAND_1328 = {1{`RANDOM}};
  field_stack_13_field_type_12_field_type = _RAND_1328[4:0];
  _RAND_1329 = {1{`RANDOM}};
  field_stack_13_field_type_12_sub_class_id = _RAND_1329[15:0];
  _RAND_1330 = {1{`RANDOM}};
  field_stack_13_field_type_13_is_repeated = _RAND_1330[0:0];
  _RAND_1331 = {1{`RANDOM}};
  field_stack_13_field_type_13_field_type = _RAND_1331[4:0];
  _RAND_1332 = {1{`RANDOM}};
  field_stack_13_field_type_13_sub_class_id = _RAND_1332[15:0];
  _RAND_1333 = {1{`RANDOM}};
  field_stack_13_field_type_14_is_repeated = _RAND_1333[0:0];
  _RAND_1334 = {1{`RANDOM}};
  field_stack_13_field_type_14_field_type = _RAND_1334[4:0];
  _RAND_1335 = {1{`RANDOM}};
  field_stack_13_field_type_14_sub_class_id = _RAND_1335[15:0];
  _RAND_1336 = {1{`RANDOM}};
  field_stack_13_field_type_15_is_repeated = _RAND_1336[0:0];
  _RAND_1337 = {1{`RANDOM}};
  field_stack_13_field_type_15_field_type = _RAND_1337[4:0];
  _RAND_1338 = {1{`RANDOM}};
  field_stack_13_field_type_15_sub_class_id = _RAND_1338[15:0];
  _RAND_1339 = {1{`RANDOM}};
  field_stack_13_field_type_16_is_repeated = _RAND_1339[0:0];
  _RAND_1340 = {1{`RANDOM}};
  field_stack_13_field_type_16_field_type = _RAND_1340[4:0];
  _RAND_1341 = {1{`RANDOM}};
  field_stack_13_field_type_16_sub_class_id = _RAND_1341[15:0];
  _RAND_1342 = {1{`RANDOM}};
  field_stack_13_field_type_17_is_repeated = _RAND_1342[0:0];
  _RAND_1343 = {1{`RANDOM}};
  field_stack_13_field_type_17_field_type = _RAND_1343[4:0];
  _RAND_1344 = {1{`RANDOM}};
  field_stack_13_field_type_17_sub_class_id = _RAND_1344[15:0];
  _RAND_1345 = {1{`RANDOM}};
  field_stack_13_field_type_18_is_repeated = _RAND_1345[0:0];
  _RAND_1346 = {1{`RANDOM}};
  field_stack_13_field_type_18_field_type = _RAND_1346[4:0];
  _RAND_1347 = {1{`RANDOM}};
  field_stack_13_field_type_18_sub_class_id = _RAND_1347[15:0];
  _RAND_1348 = {1{`RANDOM}};
  field_stack_13_field_type_19_is_repeated = _RAND_1348[0:0];
  _RAND_1349 = {1{`RANDOM}};
  field_stack_13_field_type_19_field_type = _RAND_1349[4:0];
  _RAND_1350 = {1{`RANDOM}};
  field_stack_13_field_type_19_sub_class_id = _RAND_1350[15:0];
  _RAND_1351 = {1{`RANDOM}};
  field_stack_13_field_type_20_is_repeated = _RAND_1351[0:0];
  _RAND_1352 = {1{`RANDOM}};
  field_stack_13_field_type_20_field_type = _RAND_1352[4:0];
  _RAND_1353 = {1{`RANDOM}};
  field_stack_13_field_type_20_sub_class_id = _RAND_1353[15:0];
  _RAND_1354 = {1{`RANDOM}};
  field_stack_13_field_type_21_is_repeated = _RAND_1354[0:0];
  _RAND_1355 = {1{`RANDOM}};
  field_stack_13_field_type_21_field_type = _RAND_1355[4:0];
  _RAND_1356 = {1{`RANDOM}};
  field_stack_13_field_type_21_sub_class_id = _RAND_1356[15:0];
  _RAND_1357 = {1{`RANDOM}};
  field_stack_13_field_type_22_is_repeated = _RAND_1357[0:0];
  _RAND_1358 = {1{`RANDOM}};
  field_stack_13_field_type_22_field_type = _RAND_1358[4:0];
  _RAND_1359 = {1{`RANDOM}};
  field_stack_13_field_type_22_sub_class_id = _RAND_1359[15:0];
  _RAND_1360 = {1{`RANDOM}};
  field_stack_13_field_type_23_is_repeated = _RAND_1360[0:0];
  _RAND_1361 = {1{`RANDOM}};
  field_stack_13_field_type_23_field_type = _RAND_1361[4:0];
  _RAND_1362 = {1{`RANDOM}};
  field_stack_13_field_type_23_sub_class_id = _RAND_1362[15:0];
  _RAND_1363 = {1{`RANDOM}};
  field_stack_13_field_type_24_is_repeated = _RAND_1363[0:0];
  _RAND_1364 = {1{`RANDOM}};
  field_stack_13_field_type_24_field_type = _RAND_1364[4:0];
  _RAND_1365 = {1{`RANDOM}};
  field_stack_13_field_type_24_sub_class_id = _RAND_1365[15:0];
  _RAND_1366 = {1{`RANDOM}};
  field_stack_13_field_type_25_is_repeated = _RAND_1366[0:0];
  _RAND_1367 = {1{`RANDOM}};
  field_stack_13_field_type_25_field_type = _RAND_1367[4:0];
  _RAND_1368 = {1{`RANDOM}};
  field_stack_13_field_type_25_sub_class_id = _RAND_1368[15:0];
  _RAND_1369 = {1{`RANDOM}};
  field_stack_13_field_type_26_is_repeated = _RAND_1369[0:0];
  _RAND_1370 = {1{`RANDOM}};
  field_stack_13_field_type_26_field_type = _RAND_1370[4:0];
  _RAND_1371 = {1{`RANDOM}};
  field_stack_13_field_type_26_sub_class_id = _RAND_1371[15:0];
  _RAND_1372 = {1{`RANDOM}};
  field_stack_13_field_type_27_is_repeated = _RAND_1372[0:0];
  _RAND_1373 = {1{`RANDOM}};
  field_stack_13_field_type_27_field_type = _RAND_1373[4:0];
  _RAND_1374 = {1{`RANDOM}};
  field_stack_13_field_type_27_sub_class_id = _RAND_1374[15:0];
  _RAND_1375 = {1{`RANDOM}};
  field_stack_13_field_type_28_is_repeated = _RAND_1375[0:0];
  _RAND_1376 = {1{`RANDOM}};
  field_stack_13_field_type_28_field_type = _RAND_1376[4:0];
  _RAND_1377 = {1{`RANDOM}};
  field_stack_13_field_type_28_sub_class_id = _RAND_1377[15:0];
  _RAND_1378 = {1{`RANDOM}};
  field_stack_13_field_type_29_is_repeated = _RAND_1378[0:0];
  _RAND_1379 = {1{`RANDOM}};
  field_stack_13_field_type_29_field_type = _RAND_1379[4:0];
  _RAND_1380 = {1{`RANDOM}};
  field_stack_13_field_type_29_sub_class_id = _RAND_1380[15:0];
  _RAND_1381 = {1{`RANDOM}};
  field_stack_13_field_type_30_is_repeated = _RAND_1381[0:0];
  _RAND_1382 = {1{`RANDOM}};
  field_stack_13_field_type_30_field_type = _RAND_1382[4:0];
  _RAND_1383 = {1{`RANDOM}};
  field_stack_13_field_type_30_sub_class_id = _RAND_1383[15:0];
  _RAND_1384 = {1{`RANDOM}};
  field_stack_13_field_type_31_is_repeated = _RAND_1384[0:0];
  _RAND_1385 = {1{`RANDOM}};
  field_stack_13_field_type_31_field_type = _RAND_1385[4:0];
  _RAND_1386 = {1{`RANDOM}};
  field_stack_13_field_type_31_sub_class_id = _RAND_1386[15:0];
  _RAND_1387 = {1{`RANDOM}};
  field_stack_13_field_type_32_is_repeated = _RAND_1387[0:0];
  _RAND_1388 = {1{`RANDOM}};
  field_stack_13_field_type_32_field_type = _RAND_1388[4:0];
  _RAND_1389 = {1{`RANDOM}};
  field_stack_13_field_type_32_sub_class_id = _RAND_1389[15:0];
  _RAND_1390 = {1{`RANDOM}};
  field_stack_14_field_type_0_is_repeated = _RAND_1390[0:0];
  _RAND_1391 = {1{`RANDOM}};
  field_stack_14_field_type_0_field_type = _RAND_1391[4:0];
  _RAND_1392 = {1{`RANDOM}};
  field_stack_14_field_type_0_sub_class_id = _RAND_1392[15:0];
  _RAND_1393 = {1{`RANDOM}};
  field_stack_14_field_type_1_is_repeated = _RAND_1393[0:0];
  _RAND_1394 = {1{`RANDOM}};
  field_stack_14_field_type_1_field_type = _RAND_1394[4:0];
  _RAND_1395 = {1{`RANDOM}};
  field_stack_14_field_type_1_sub_class_id = _RAND_1395[15:0];
  _RAND_1396 = {1{`RANDOM}};
  field_stack_14_field_type_2_is_repeated = _RAND_1396[0:0];
  _RAND_1397 = {1{`RANDOM}};
  field_stack_14_field_type_2_field_type = _RAND_1397[4:0];
  _RAND_1398 = {1{`RANDOM}};
  field_stack_14_field_type_2_sub_class_id = _RAND_1398[15:0];
  _RAND_1399 = {1{`RANDOM}};
  field_stack_14_field_type_3_is_repeated = _RAND_1399[0:0];
  _RAND_1400 = {1{`RANDOM}};
  field_stack_14_field_type_3_field_type = _RAND_1400[4:0];
  _RAND_1401 = {1{`RANDOM}};
  field_stack_14_field_type_3_sub_class_id = _RAND_1401[15:0];
  _RAND_1402 = {1{`RANDOM}};
  field_stack_14_field_type_4_is_repeated = _RAND_1402[0:0];
  _RAND_1403 = {1{`RANDOM}};
  field_stack_14_field_type_4_field_type = _RAND_1403[4:0];
  _RAND_1404 = {1{`RANDOM}};
  field_stack_14_field_type_4_sub_class_id = _RAND_1404[15:0];
  _RAND_1405 = {1{`RANDOM}};
  field_stack_14_field_type_5_is_repeated = _RAND_1405[0:0];
  _RAND_1406 = {1{`RANDOM}};
  field_stack_14_field_type_5_field_type = _RAND_1406[4:0];
  _RAND_1407 = {1{`RANDOM}};
  field_stack_14_field_type_5_sub_class_id = _RAND_1407[15:0];
  _RAND_1408 = {1{`RANDOM}};
  field_stack_14_field_type_6_is_repeated = _RAND_1408[0:0];
  _RAND_1409 = {1{`RANDOM}};
  field_stack_14_field_type_6_field_type = _RAND_1409[4:0];
  _RAND_1410 = {1{`RANDOM}};
  field_stack_14_field_type_6_sub_class_id = _RAND_1410[15:0];
  _RAND_1411 = {1{`RANDOM}};
  field_stack_14_field_type_7_is_repeated = _RAND_1411[0:0];
  _RAND_1412 = {1{`RANDOM}};
  field_stack_14_field_type_7_field_type = _RAND_1412[4:0];
  _RAND_1413 = {1{`RANDOM}};
  field_stack_14_field_type_7_sub_class_id = _RAND_1413[15:0];
  _RAND_1414 = {1{`RANDOM}};
  field_stack_14_field_type_8_is_repeated = _RAND_1414[0:0];
  _RAND_1415 = {1{`RANDOM}};
  field_stack_14_field_type_8_field_type = _RAND_1415[4:0];
  _RAND_1416 = {1{`RANDOM}};
  field_stack_14_field_type_8_sub_class_id = _RAND_1416[15:0];
  _RAND_1417 = {1{`RANDOM}};
  field_stack_14_field_type_9_is_repeated = _RAND_1417[0:0];
  _RAND_1418 = {1{`RANDOM}};
  field_stack_14_field_type_9_field_type = _RAND_1418[4:0];
  _RAND_1419 = {1{`RANDOM}};
  field_stack_14_field_type_9_sub_class_id = _RAND_1419[15:0];
  _RAND_1420 = {1{`RANDOM}};
  field_stack_14_field_type_10_is_repeated = _RAND_1420[0:0];
  _RAND_1421 = {1{`RANDOM}};
  field_stack_14_field_type_10_field_type = _RAND_1421[4:0];
  _RAND_1422 = {1{`RANDOM}};
  field_stack_14_field_type_10_sub_class_id = _RAND_1422[15:0];
  _RAND_1423 = {1{`RANDOM}};
  field_stack_14_field_type_11_is_repeated = _RAND_1423[0:0];
  _RAND_1424 = {1{`RANDOM}};
  field_stack_14_field_type_11_field_type = _RAND_1424[4:0];
  _RAND_1425 = {1{`RANDOM}};
  field_stack_14_field_type_11_sub_class_id = _RAND_1425[15:0];
  _RAND_1426 = {1{`RANDOM}};
  field_stack_14_field_type_12_is_repeated = _RAND_1426[0:0];
  _RAND_1427 = {1{`RANDOM}};
  field_stack_14_field_type_12_field_type = _RAND_1427[4:0];
  _RAND_1428 = {1{`RANDOM}};
  field_stack_14_field_type_12_sub_class_id = _RAND_1428[15:0];
  _RAND_1429 = {1{`RANDOM}};
  field_stack_14_field_type_13_is_repeated = _RAND_1429[0:0];
  _RAND_1430 = {1{`RANDOM}};
  field_stack_14_field_type_13_field_type = _RAND_1430[4:0];
  _RAND_1431 = {1{`RANDOM}};
  field_stack_14_field_type_13_sub_class_id = _RAND_1431[15:0];
  _RAND_1432 = {1{`RANDOM}};
  field_stack_14_field_type_14_is_repeated = _RAND_1432[0:0];
  _RAND_1433 = {1{`RANDOM}};
  field_stack_14_field_type_14_field_type = _RAND_1433[4:0];
  _RAND_1434 = {1{`RANDOM}};
  field_stack_14_field_type_14_sub_class_id = _RAND_1434[15:0];
  _RAND_1435 = {1{`RANDOM}};
  field_stack_14_field_type_15_is_repeated = _RAND_1435[0:0];
  _RAND_1436 = {1{`RANDOM}};
  field_stack_14_field_type_15_field_type = _RAND_1436[4:0];
  _RAND_1437 = {1{`RANDOM}};
  field_stack_14_field_type_15_sub_class_id = _RAND_1437[15:0];
  _RAND_1438 = {1{`RANDOM}};
  field_stack_14_field_type_16_is_repeated = _RAND_1438[0:0];
  _RAND_1439 = {1{`RANDOM}};
  field_stack_14_field_type_16_field_type = _RAND_1439[4:0];
  _RAND_1440 = {1{`RANDOM}};
  field_stack_14_field_type_16_sub_class_id = _RAND_1440[15:0];
  _RAND_1441 = {1{`RANDOM}};
  field_stack_14_field_type_17_is_repeated = _RAND_1441[0:0];
  _RAND_1442 = {1{`RANDOM}};
  field_stack_14_field_type_17_field_type = _RAND_1442[4:0];
  _RAND_1443 = {1{`RANDOM}};
  field_stack_14_field_type_17_sub_class_id = _RAND_1443[15:0];
  _RAND_1444 = {1{`RANDOM}};
  field_stack_14_field_type_18_is_repeated = _RAND_1444[0:0];
  _RAND_1445 = {1{`RANDOM}};
  field_stack_14_field_type_18_field_type = _RAND_1445[4:0];
  _RAND_1446 = {1{`RANDOM}};
  field_stack_14_field_type_18_sub_class_id = _RAND_1446[15:0];
  _RAND_1447 = {1{`RANDOM}};
  field_stack_14_field_type_19_is_repeated = _RAND_1447[0:0];
  _RAND_1448 = {1{`RANDOM}};
  field_stack_14_field_type_19_field_type = _RAND_1448[4:0];
  _RAND_1449 = {1{`RANDOM}};
  field_stack_14_field_type_19_sub_class_id = _RAND_1449[15:0];
  _RAND_1450 = {1{`RANDOM}};
  field_stack_14_field_type_20_is_repeated = _RAND_1450[0:0];
  _RAND_1451 = {1{`RANDOM}};
  field_stack_14_field_type_20_field_type = _RAND_1451[4:0];
  _RAND_1452 = {1{`RANDOM}};
  field_stack_14_field_type_20_sub_class_id = _RAND_1452[15:0];
  _RAND_1453 = {1{`RANDOM}};
  field_stack_14_field_type_21_is_repeated = _RAND_1453[0:0];
  _RAND_1454 = {1{`RANDOM}};
  field_stack_14_field_type_21_field_type = _RAND_1454[4:0];
  _RAND_1455 = {1{`RANDOM}};
  field_stack_14_field_type_21_sub_class_id = _RAND_1455[15:0];
  _RAND_1456 = {1{`RANDOM}};
  field_stack_14_field_type_22_is_repeated = _RAND_1456[0:0];
  _RAND_1457 = {1{`RANDOM}};
  field_stack_14_field_type_22_field_type = _RAND_1457[4:0];
  _RAND_1458 = {1{`RANDOM}};
  field_stack_14_field_type_22_sub_class_id = _RAND_1458[15:0];
  _RAND_1459 = {1{`RANDOM}};
  field_stack_14_field_type_23_is_repeated = _RAND_1459[0:0];
  _RAND_1460 = {1{`RANDOM}};
  field_stack_14_field_type_23_field_type = _RAND_1460[4:0];
  _RAND_1461 = {1{`RANDOM}};
  field_stack_14_field_type_23_sub_class_id = _RAND_1461[15:0];
  _RAND_1462 = {1{`RANDOM}};
  field_stack_14_field_type_24_is_repeated = _RAND_1462[0:0];
  _RAND_1463 = {1{`RANDOM}};
  field_stack_14_field_type_24_field_type = _RAND_1463[4:0];
  _RAND_1464 = {1{`RANDOM}};
  field_stack_14_field_type_24_sub_class_id = _RAND_1464[15:0];
  _RAND_1465 = {1{`RANDOM}};
  field_stack_14_field_type_25_is_repeated = _RAND_1465[0:0];
  _RAND_1466 = {1{`RANDOM}};
  field_stack_14_field_type_25_field_type = _RAND_1466[4:0];
  _RAND_1467 = {1{`RANDOM}};
  field_stack_14_field_type_25_sub_class_id = _RAND_1467[15:0];
  _RAND_1468 = {1{`RANDOM}};
  field_stack_14_field_type_26_is_repeated = _RAND_1468[0:0];
  _RAND_1469 = {1{`RANDOM}};
  field_stack_14_field_type_26_field_type = _RAND_1469[4:0];
  _RAND_1470 = {1{`RANDOM}};
  field_stack_14_field_type_26_sub_class_id = _RAND_1470[15:0];
  _RAND_1471 = {1{`RANDOM}};
  field_stack_14_field_type_27_is_repeated = _RAND_1471[0:0];
  _RAND_1472 = {1{`RANDOM}};
  field_stack_14_field_type_27_field_type = _RAND_1472[4:0];
  _RAND_1473 = {1{`RANDOM}};
  field_stack_14_field_type_27_sub_class_id = _RAND_1473[15:0];
  _RAND_1474 = {1{`RANDOM}};
  field_stack_14_field_type_28_is_repeated = _RAND_1474[0:0];
  _RAND_1475 = {1{`RANDOM}};
  field_stack_14_field_type_28_field_type = _RAND_1475[4:0];
  _RAND_1476 = {1{`RANDOM}};
  field_stack_14_field_type_28_sub_class_id = _RAND_1476[15:0];
  _RAND_1477 = {1{`RANDOM}};
  field_stack_14_field_type_29_is_repeated = _RAND_1477[0:0];
  _RAND_1478 = {1{`RANDOM}};
  field_stack_14_field_type_29_field_type = _RAND_1478[4:0];
  _RAND_1479 = {1{`RANDOM}};
  field_stack_14_field_type_29_sub_class_id = _RAND_1479[15:0];
  _RAND_1480 = {1{`RANDOM}};
  field_stack_14_field_type_30_is_repeated = _RAND_1480[0:0];
  _RAND_1481 = {1{`RANDOM}};
  field_stack_14_field_type_30_field_type = _RAND_1481[4:0];
  _RAND_1482 = {1{`RANDOM}};
  field_stack_14_field_type_30_sub_class_id = _RAND_1482[15:0];
  _RAND_1483 = {1{`RANDOM}};
  field_stack_14_field_type_31_is_repeated = _RAND_1483[0:0];
  _RAND_1484 = {1{`RANDOM}};
  field_stack_14_field_type_31_field_type = _RAND_1484[4:0];
  _RAND_1485 = {1{`RANDOM}};
  field_stack_14_field_type_31_sub_class_id = _RAND_1485[15:0];
  _RAND_1486 = {1{`RANDOM}};
  field_stack_14_field_type_32_is_repeated = _RAND_1486[0:0];
  _RAND_1487 = {1{`RANDOM}};
  field_stack_14_field_type_32_field_type = _RAND_1487[4:0];
  _RAND_1488 = {1{`RANDOM}};
  field_stack_14_field_type_32_sub_class_id = _RAND_1488[15:0];
  _RAND_1489 = {1{`RANDOM}};
  field_num_0 = _RAND_1489[5:0];
  _RAND_1490 = {1{`RANDOM}};
  field_num_1 = _RAND_1490[5:0];
  _RAND_1491 = {1{`RANDOM}};
  field_num_2 = _RAND_1491[5:0];
  _RAND_1492 = {1{`RANDOM}};
  field_num_3 = _RAND_1492[5:0];
  _RAND_1493 = {1{`RANDOM}};
  field_num_4 = _RAND_1493[5:0];
  _RAND_1494 = {1{`RANDOM}};
  field_num_5 = _RAND_1494[5:0];
  _RAND_1495 = {1{`RANDOM}};
  field_num_6 = _RAND_1495[5:0];
  _RAND_1496 = {1{`RANDOM}};
  field_num_7 = _RAND_1496[5:0];
  _RAND_1497 = {1{`RANDOM}};
  field_num_8 = _RAND_1497[5:0];
  _RAND_1498 = {1{`RANDOM}};
  field_num_9 = _RAND_1498[5:0];
  _RAND_1499 = {1{`RANDOM}};
  field_num_10 = _RAND_1499[5:0];
  _RAND_1500 = {1{`RANDOM}};
  field_num_11 = _RAND_1500[5:0];
  _RAND_1501 = {1{`RANDOM}};
  field_num_12 = _RAND_1501[5:0];
  _RAND_1502 = {1{`RANDOM}};
  field_num_13 = _RAND_1502[5:0];
  _RAND_1503 = {1{`RANDOM}};
  field_num_14 = _RAND_1503[5:0];
  _RAND_1504 = {1{`RANDOM}};
  field_num_15 = _RAND_1504[5:0];
  _RAND_1505 = {2{`RANDOM}};
  host_base_addr = _RAND_1505[63:0];
  _RAND_1506 = {1{`RANDOM}};
  current_field_num = _RAND_1506[5:0];
  _RAND_1507 = {1{`RANDOM}};
  c_sub_metadata_is_repeated = _RAND_1507[0:0];
  _RAND_1508 = {1{`RANDOM}};
  c_sub_metadata_field_type = _RAND_1508[4:0];
  _RAND_1509 = {1{`RANDOM}};
  c_sub_metadata_sub_class_id = _RAND_1509[15:0];
  _RAND_1510 = {1{`RANDOM}};
  repeat_num = _RAND_1510[7:0];
  _RAND_1511 = {1{`RANDOM}};
  stack_num = _RAND_1511[3:0];
  _RAND_1512 = {1{`RANDOM}};
  current_field_length = _RAND_1512[31:0];
  _RAND_1513 = {1{`RANDOM}};
  state = _RAND_1513[4:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Queue_6(
  input        clock,
  input        reset,
  output       io_enq_ready,
  input        io_enq_valid,
  input  [9:0] io_enq_bits_class_id,
  input        io_deq_ready,
  output       io_deq_valid,
  output [9:0] io_deq_bits_class_id
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
`endif // RANDOMIZE_REG_INIT
  reg [9:0] ram_class_id [0:7]; // @[Decoupled.scala 218:16]
  wire [9:0] ram_class_id_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16]
  wire [2:0] ram_class_id_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16]
  wire [9:0] ram_class_id_MPORT_data; // @[Decoupled.scala 218:16]
  wire [2:0] ram_class_id_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_class_id_MPORT_mask; // @[Decoupled.scala 218:16]
  wire  ram_class_id_MPORT_en; // @[Decoupled.scala 218:16]
  reg [2:0] enq_ptr_value; // @[Counter.scala 60:40]
  reg [2:0] deq_ptr_value; // @[Counter.scala 60:40]
  reg  maybe_full; // @[Decoupled.scala 221:27]
  wire  ptr_match = enq_ptr_value == deq_ptr_value; // @[Decoupled.scala 223:33]
  wire  empty = ptr_match & ~maybe_full; // @[Decoupled.scala 224:25]
  wire  full = ptr_match & maybe_full; // @[Decoupled.scala 225:24]
  wire  do_enq = io_enq_ready & io_enq_valid; // @[Decoupled.scala 40:37]
  wire  do_deq = io_deq_ready & io_deq_valid; // @[Decoupled.scala 40:37]
  wire [2:0] _value_T_1 = enq_ptr_value + 3'h1; // @[Counter.scala 76:24]
  wire [2:0] _value_T_3 = deq_ptr_value + 3'h1; // @[Counter.scala 76:24]
  assign ram_class_id_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_class_id_io_deq_bits_MPORT_data = ram_class_id[ram_class_id_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  assign ram_class_id_MPORT_data = io_enq_bits_class_id;
  assign ram_class_id_MPORT_addr = enq_ptr_value;
  assign ram_class_id_MPORT_mask = 1'h1;
  assign ram_class_id_MPORT_en = io_enq_ready & io_enq_valid;
  assign io_enq_ready = ~full; // @[Decoupled.scala 241:19]
  assign io_deq_valid = ~empty; // @[Decoupled.scala 240:19]
  assign io_deq_bits_class_id = ram_class_id_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15]
  always @(posedge clock) begin
    if(ram_class_id_MPORT_en & ram_class_id_MPORT_mask) begin
      ram_class_id[ram_class_id_MPORT_addr] <= ram_class_id_MPORT_data; // @[Decoupled.scala 218:16]
    end
    if (reset) begin // @[Counter.scala 60:40]
      enq_ptr_value <= 3'h0; // @[Counter.scala 60:40]
    end else if (do_enq) begin // @[Decoupled.scala 229:17]
      enq_ptr_value <= _value_T_1; // @[Counter.scala 76:15]
    end
    if (reset) begin // @[Counter.scala 60:40]
      deq_ptr_value <= 3'h0; // @[Counter.scala 60:40]
    end else if (do_deq) begin // @[Decoupled.scala 233:17]
      deq_ptr_value <= _value_T_3; // @[Counter.scala 76:15]
    end
    if (reset) begin // @[Decoupled.scala 221:27]
      maybe_full <= 1'h0; // @[Decoupled.scala 221:27]
    end else if (do_enq != do_deq) begin // @[Decoupled.scala 236:28]
      maybe_full <= do_enq; // @[Decoupled.scala 237:16]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 8; initvar = initvar+1)
    ram_class_id[initvar] = _RAND_0[9:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  enq_ptr_value = _RAND_1[2:0];
  _RAND_2 = {1{`RANDOM}};
  deq_ptr_value = _RAND_2[2:0];
  _RAND_3 = {1{`RANDOM}};
  maybe_full = _RAND_3[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module XQueue_4(
  input        clock,
  input        reset,
  output       io_in_ready,
  input        io_in_valid,
  input  [9:0] io_in_bits_class_id,
  input        io_out_ready,
  output       io_out_valid,
  output [9:0] io_out_bits_class_id
);
  wire  q_clock; // @[XQueue.scala 85:39]
  wire  q_reset; // @[XQueue.scala 85:39]
  wire  q_io_enq_ready; // @[XQueue.scala 85:39]
  wire  q_io_enq_valid; // @[XQueue.scala 85:39]
  wire [9:0] q_io_enq_bits_class_id; // @[XQueue.scala 85:39]
  wire  q_io_deq_ready; // @[XQueue.scala 85:39]
  wire  q_io_deq_valid; // @[XQueue.scala 85:39]
  wire [9:0] q_io_deq_bits_class_id; // @[XQueue.scala 85:39]
  Queue_6 q ( // @[XQueue.scala 85:39]
    .clock(q_clock),
    .reset(q_reset),
    .io_enq_ready(q_io_enq_ready),
    .io_enq_valid(q_io_enq_valid),
    .io_enq_bits_class_id(q_io_enq_bits_class_id),
    .io_deq_ready(q_io_deq_ready),
    .io_deq_valid(q_io_deq_valid),
    .io_deq_bits_class_id(q_io_deq_bits_class_id)
  );
  assign io_in_ready = q_io_enq_ready; // @[XQueue.scala 87:34]
  assign io_out_valid = q_io_deq_valid; // @[XQueue.scala 88:34]
  assign io_out_bits_class_id = q_io_deq_bits_class_id; // @[XQueue.scala 88:34]
  assign q_clock = clock;
  assign q_reset = reset;
  assign q_io_enq_valid = io_in_valid; // @[XQueue.scala 87:34]
  assign q_io_enq_bits_class_id = io_in_bits_class_id; // @[XQueue.scala 87:34]
  assign q_io_deq_ready = io_out_ready; // @[XQueue.scala 88:34]
endmodule
module XRam_1(
  input         clock,
  input         reset,
  input  [9:0]  io_addr_a,
  input  [9:0]  io_addr_b,
  input         io_wr_en_a,
  input  [15:0] io_data_in_a_class_length,
  input  [7:0]  io_data_in_a_max_field_num,
  input         io_data_in_a_field_type_0_is_repeated,
  input  [4:0]  io_data_in_a_field_type_0_field_type,
  input  [15:0] io_data_in_a_field_type_0_sub_class_id,
  input         io_data_in_a_field_type_0_is_host,
  input         io_data_in_a_field_type_1_is_repeated,
  input  [4:0]  io_data_in_a_field_type_1_field_type,
  input  [15:0] io_data_in_a_field_type_1_sub_class_id,
  input         io_data_in_a_field_type_1_is_host,
  input         io_data_in_a_field_type_2_is_repeated,
  input  [4:0]  io_data_in_a_field_type_2_field_type,
  input  [15:0] io_data_in_a_field_type_2_sub_class_id,
  input         io_data_in_a_field_type_2_is_host,
  input         io_data_in_a_field_type_3_is_repeated,
  input  [4:0]  io_data_in_a_field_type_3_field_type,
  input  [15:0] io_data_in_a_field_type_3_sub_class_id,
  input         io_data_in_a_field_type_3_is_host,
  input         io_data_in_a_field_type_4_is_repeated,
  input  [4:0]  io_data_in_a_field_type_4_field_type,
  input  [15:0] io_data_in_a_field_type_4_sub_class_id,
  input         io_data_in_a_field_type_4_is_host,
  input         io_data_in_a_field_type_5_is_repeated,
  input  [4:0]  io_data_in_a_field_type_5_field_type,
  input  [15:0] io_data_in_a_field_type_5_sub_class_id,
  input         io_data_in_a_field_type_5_is_host,
  input         io_data_in_a_field_type_6_is_repeated,
  input  [4:0]  io_data_in_a_field_type_6_field_type,
  input  [15:0] io_data_in_a_field_type_6_sub_class_id,
  input         io_data_in_a_field_type_6_is_host,
  input         io_data_in_a_field_type_7_is_repeated,
  input  [4:0]  io_data_in_a_field_type_7_field_type,
  input  [15:0] io_data_in_a_field_type_7_sub_class_id,
  input         io_data_in_a_field_type_7_is_host,
  input         io_data_in_a_field_type_8_is_repeated,
  input  [4:0]  io_data_in_a_field_type_8_field_type,
  input  [15:0] io_data_in_a_field_type_8_sub_class_id,
  input         io_data_in_a_field_type_8_is_host,
  input         io_data_in_a_field_type_9_is_repeated,
  input  [4:0]  io_data_in_a_field_type_9_field_type,
  input  [15:0] io_data_in_a_field_type_9_sub_class_id,
  input         io_data_in_a_field_type_9_is_host,
  input         io_data_in_a_field_type_10_is_repeated,
  input  [4:0]  io_data_in_a_field_type_10_field_type,
  input  [15:0] io_data_in_a_field_type_10_sub_class_id,
  input         io_data_in_a_field_type_10_is_host,
  input         io_data_in_a_field_type_11_is_repeated,
  input  [4:0]  io_data_in_a_field_type_11_field_type,
  input  [15:0] io_data_in_a_field_type_11_sub_class_id,
  input         io_data_in_a_field_type_11_is_host,
  input         io_data_in_a_field_type_12_is_repeated,
  input  [4:0]  io_data_in_a_field_type_12_field_type,
  input  [15:0] io_data_in_a_field_type_12_sub_class_id,
  input         io_data_in_a_field_type_12_is_host,
  input         io_data_in_a_field_type_13_is_repeated,
  input  [4:0]  io_data_in_a_field_type_13_field_type,
  input  [15:0] io_data_in_a_field_type_13_sub_class_id,
  input         io_data_in_a_field_type_13_is_host,
  input         io_data_in_a_field_type_14_is_repeated,
  input  [4:0]  io_data_in_a_field_type_14_field_type,
  input  [15:0] io_data_in_a_field_type_14_sub_class_id,
  input         io_data_in_a_field_type_14_is_host,
  input         io_data_in_a_field_type_15_is_repeated,
  input  [4:0]  io_data_in_a_field_type_15_field_type,
  input  [15:0] io_data_in_a_field_type_15_sub_class_id,
  input         io_data_in_a_field_type_15_is_host,
  input         io_data_in_a_field_type_16_is_repeated,
  input  [4:0]  io_data_in_a_field_type_16_field_type,
  input  [15:0] io_data_in_a_field_type_16_sub_class_id,
  input         io_data_in_a_field_type_16_is_host,
  input         io_data_in_a_field_type_17_is_repeated,
  input  [4:0]  io_data_in_a_field_type_17_field_type,
  input  [15:0] io_data_in_a_field_type_17_sub_class_id,
  input         io_data_in_a_field_type_17_is_host,
  input         io_data_in_a_field_type_18_is_repeated,
  input  [4:0]  io_data_in_a_field_type_18_field_type,
  input  [15:0] io_data_in_a_field_type_18_sub_class_id,
  input         io_data_in_a_field_type_18_is_host,
  input         io_data_in_a_field_type_19_is_repeated,
  input  [4:0]  io_data_in_a_field_type_19_field_type,
  input  [15:0] io_data_in_a_field_type_19_sub_class_id,
  input         io_data_in_a_field_type_19_is_host,
  input         io_data_in_a_field_type_20_is_repeated,
  input  [4:0]  io_data_in_a_field_type_20_field_type,
  input  [15:0] io_data_in_a_field_type_20_sub_class_id,
  input         io_data_in_a_field_type_20_is_host,
  input         io_data_in_a_field_type_21_is_repeated,
  input  [4:0]  io_data_in_a_field_type_21_field_type,
  input  [15:0] io_data_in_a_field_type_21_sub_class_id,
  input         io_data_in_a_field_type_21_is_host,
  input         io_data_in_a_field_type_22_is_repeated,
  input  [4:0]  io_data_in_a_field_type_22_field_type,
  input  [15:0] io_data_in_a_field_type_22_sub_class_id,
  input         io_data_in_a_field_type_22_is_host,
  input         io_data_in_a_field_type_23_is_repeated,
  input  [4:0]  io_data_in_a_field_type_23_field_type,
  input  [15:0] io_data_in_a_field_type_23_sub_class_id,
  input         io_data_in_a_field_type_23_is_host,
  input         io_data_in_a_field_type_24_is_repeated,
  input  [4:0]  io_data_in_a_field_type_24_field_type,
  input  [15:0] io_data_in_a_field_type_24_sub_class_id,
  input         io_data_in_a_field_type_24_is_host,
  input         io_data_in_a_field_type_25_is_repeated,
  input  [4:0]  io_data_in_a_field_type_25_field_type,
  input  [15:0] io_data_in_a_field_type_25_sub_class_id,
  input         io_data_in_a_field_type_25_is_host,
  input         io_data_in_a_field_type_26_is_repeated,
  input  [4:0]  io_data_in_a_field_type_26_field_type,
  input  [15:0] io_data_in_a_field_type_26_sub_class_id,
  input         io_data_in_a_field_type_26_is_host,
  input         io_data_in_a_field_type_27_is_repeated,
  input  [4:0]  io_data_in_a_field_type_27_field_type,
  input  [15:0] io_data_in_a_field_type_27_sub_class_id,
  input         io_data_in_a_field_type_27_is_host,
  input         io_data_in_a_field_type_28_is_repeated,
  input  [4:0]  io_data_in_a_field_type_28_field_type,
  input  [15:0] io_data_in_a_field_type_28_sub_class_id,
  input         io_data_in_a_field_type_28_is_host,
  input         io_data_in_a_field_type_29_is_repeated,
  input  [4:0]  io_data_in_a_field_type_29_field_type,
  input  [15:0] io_data_in_a_field_type_29_sub_class_id,
  input         io_data_in_a_field_type_29_is_host,
  input         io_data_in_a_field_type_30_is_repeated,
  input  [4:0]  io_data_in_a_field_type_30_field_type,
  input  [15:0] io_data_in_a_field_type_30_sub_class_id,
  input         io_data_in_a_field_type_30_is_host,
  input         io_data_in_a_field_type_31_is_repeated,
  input  [4:0]  io_data_in_a_field_type_31_field_type,
  input  [15:0] io_data_in_a_field_type_31_sub_class_id,
  input         io_data_in_a_field_type_31_is_host,
  input         io_data_in_a_field_type_32_is_repeated,
  input  [4:0]  io_data_in_a_field_type_32_field_type,
  input  [15:0] io_data_in_a_field_type_32_sub_class_id,
  input         io_data_in_a_field_type_32_is_host,
  output [7:0]  io_data_out_b_max_field_num,
  output        io_data_out_b_field_type_0_is_repeated,
  output [4:0]  io_data_out_b_field_type_0_field_type,
  output [15:0] io_data_out_b_field_type_0_sub_class_id,
  output        io_data_out_b_field_type_1_is_repeated,
  output [4:0]  io_data_out_b_field_type_1_field_type,
  output [15:0] io_data_out_b_field_type_1_sub_class_id,
  output        io_data_out_b_field_type_2_is_repeated,
  output [4:0]  io_data_out_b_field_type_2_field_type,
  output [15:0] io_data_out_b_field_type_2_sub_class_id,
  output        io_data_out_b_field_type_3_is_repeated,
  output [4:0]  io_data_out_b_field_type_3_field_type,
  output [15:0] io_data_out_b_field_type_3_sub_class_id,
  output        io_data_out_b_field_type_4_is_repeated,
  output [4:0]  io_data_out_b_field_type_4_field_type,
  output [15:0] io_data_out_b_field_type_4_sub_class_id,
  output        io_data_out_b_field_type_5_is_repeated,
  output [4:0]  io_data_out_b_field_type_5_field_type,
  output [15:0] io_data_out_b_field_type_5_sub_class_id,
  output        io_data_out_b_field_type_6_is_repeated,
  output [4:0]  io_data_out_b_field_type_6_field_type,
  output [15:0] io_data_out_b_field_type_6_sub_class_id,
  output        io_data_out_b_field_type_7_is_repeated,
  output [4:0]  io_data_out_b_field_type_7_field_type,
  output [15:0] io_data_out_b_field_type_7_sub_class_id,
  output        io_data_out_b_field_type_8_is_repeated,
  output [4:0]  io_data_out_b_field_type_8_field_type,
  output [15:0] io_data_out_b_field_type_8_sub_class_id,
  output        io_data_out_b_field_type_9_is_repeated,
  output [4:0]  io_data_out_b_field_type_9_field_type,
  output [15:0] io_data_out_b_field_type_9_sub_class_id,
  output        io_data_out_b_field_type_10_is_repeated,
  output [4:0]  io_data_out_b_field_type_10_field_type,
  output [15:0] io_data_out_b_field_type_10_sub_class_id,
  output        io_data_out_b_field_type_11_is_repeated,
  output [4:0]  io_data_out_b_field_type_11_field_type,
  output [15:0] io_data_out_b_field_type_11_sub_class_id,
  output        io_data_out_b_field_type_12_is_repeated,
  output [4:0]  io_data_out_b_field_type_12_field_type,
  output [15:0] io_data_out_b_field_type_12_sub_class_id,
  output        io_data_out_b_field_type_13_is_repeated,
  output [4:0]  io_data_out_b_field_type_13_field_type,
  output [15:0] io_data_out_b_field_type_13_sub_class_id,
  output        io_data_out_b_field_type_14_is_repeated,
  output [4:0]  io_data_out_b_field_type_14_field_type,
  output [15:0] io_data_out_b_field_type_14_sub_class_id,
  output        io_data_out_b_field_type_15_is_repeated,
  output [4:0]  io_data_out_b_field_type_15_field_type,
  output [15:0] io_data_out_b_field_type_15_sub_class_id,
  output        io_data_out_b_field_type_16_is_repeated,
  output [4:0]  io_data_out_b_field_type_16_field_type,
  output [15:0] io_data_out_b_field_type_16_sub_class_id,
  output        io_data_out_b_field_type_17_is_repeated,
  output [4:0]  io_data_out_b_field_type_17_field_type,
  output [15:0] io_data_out_b_field_type_17_sub_class_id,
  output        io_data_out_b_field_type_18_is_repeated,
  output [4:0]  io_data_out_b_field_type_18_field_type,
  output [15:0] io_data_out_b_field_type_18_sub_class_id,
  output        io_data_out_b_field_type_19_is_repeated,
  output [4:0]  io_data_out_b_field_type_19_field_type,
  output [15:0] io_data_out_b_field_type_19_sub_class_id,
  output        io_data_out_b_field_type_20_is_repeated,
  output [4:0]  io_data_out_b_field_type_20_field_type,
  output [15:0] io_data_out_b_field_type_20_sub_class_id,
  output        io_data_out_b_field_type_21_is_repeated,
  output [4:0]  io_data_out_b_field_type_21_field_type,
  output [15:0] io_data_out_b_field_type_21_sub_class_id,
  output        io_data_out_b_field_type_22_is_repeated,
  output [4:0]  io_data_out_b_field_type_22_field_type,
  output [15:0] io_data_out_b_field_type_22_sub_class_id,
  output        io_data_out_b_field_type_23_is_repeated,
  output [4:0]  io_data_out_b_field_type_23_field_type,
  output [15:0] io_data_out_b_field_type_23_sub_class_id,
  output        io_data_out_b_field_type_24_is_repeated,
  output [4:0]  io_data_out_b_field_type_24_field_type,
  output [15:0] io_data_out_b_field_type_24_sub_class_id,
  output        io_data_out_b_field_type_25_is_repeated,
  output [4:0]  io_data_out_b_field_type_25_field_type,
  output [15:0] io_data_out_b_field_type_25_sub_class_id,
  output        io_data_out_b_field_type_26_is_repeated,
  output [4:0]  io_data_out_b_field_type_26_field_type,
  output [15:0] io_data_out_b_field_type_26_sub_class_id,
  output        io_data_out_b_field_type_27_is_repeated,
  output [4:0]  io_data_out_b_field_type_27_field_type,
  output [15:0] io_data_out_b_field_type_27_sub_class_id,
  output        io_data_out_b_field_type_28_is_repeated,
  output [4:0]  io_data_out_b_field_type_28_field_type,
  output [15:0] io_data_out_b_field_type_28_sub_class_id,
  output        io_data_out_b_field_type_29_is_repeated,
  output [4:0]  io_data_out_b_field_type_29_field_type,
  output [15:0] io_data_out_b_field_type_29_sub_class_id,
  output        io_data_out_b_field_type_30_is_repeated,
  output [4:0]  io_data_out_b_field_type_30_field_type,
  output [15:0] io_data_out_b_field_type_30_sub_class_id,
  output        io_data_out_b_field_type_31_is_repeated,
  output [4:0]  io_data_out_b_field_type_31_field_type,
  output [15:0] io_data_out_b_field_type_31_sub_class_id,
  output        io_data_out_b_field_type_32_is_repeated,
  output [4:0]  io_data_out_b_field_type_32_field_type,
  output [15:0] io_data_out_b_field_type_32_sub_class_id
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
`endif // RANDOMIZE_REG_INIT
  wire [783:0] ram_douta; // @[XRam.scala 136:33]
  wire [783:0] ram_doutb; // @[XRam.scala 136:33]
  wire [9:0] ram_addra; // @[XRam.scala 136:33]
  wire [9:0] ram_addrb; // @[XRam.scala 136:33]
  wire  ram_clka; // @[XRam.scala 136:33]
  wire  ram_clkb; // @[XRam.scala 136:33]
  wire [783:0] ram_dina; // @[XRam.scala 136:33]
  wire [783:0] ram_dinb; // @[XRam.scala 136:33]
  wire  ram_ena; // @[XRam.scala 136:33]
  wire  ram_enb; // @[XRam.scala 136:33]
  wire  ram_injectdbiterra; // @[XRam.scala 136:33]
  wire  ram_injectdbiterrb; // @[XRam.scala 136:33]
  wire  ram_injectsbiterra; // @[XRam.scala 136:33]
  wire  ram_injectsbiterrb; // @[XRam.scala 136:33]
  wire  ram_regcea; // @[XRam.scala 136:33]
  wire  ram_regceb; // @[XRam.scala 136:33]
  wire  ram_rsta; // @[XRam.scala 136:33]
  wire  ram_rstb; // @[XRam.scala 136:33]
  wire  ram_sleep; // @[XRam.scala 136:33]
  wire [97:0] ram_wea; // @[XRam.scala 136:33]
  wire [97:0] ram_web; // @[XRam.scala 136:33]
  wire [97:0] wr_en_a = io_wr_en_a ? 98'h3ffffffffffffffffffffffff : 98'h0; // @[Bitwise.scala 72:12]
  reg  usr_rst_delay_r; // @[Reg.scala 15:16]
  reg  usr_rst_delay_r_1; // @[Reg.scala 15:16]
  reg  usr_rst_delay_r_2; // @[Reg.scala 15:16]
  reg  usr_rst_delay; // @[Reg.scala 15:16]
  reg [9:0] reset_addr; // @[XRam.scala 141:54]
  wire [9:0] _reset_addr_T_1 = reset_addr + 10'h1; // @[XRam.scala 144:70]
  reg [9:0] REG; // @[XRam.scala 159:45]
  reg [9:0] REG_1; // @[XRam.scala 159:68]
  reg  REG_2; // @[XRam.scala 159:89]
  reg [7:0] io_data_out_b_REG_max_field_num; // @[XRam.scala 160:75]
  reg  io_data_out_b_REG_field_type_0_is_repeated; // @[XRam.scala 160:75]
  reg [4:0] io_data_out_b_REG_field_type_0_field_type; // @[XRam.scala 160:75]
  reg [15:0] io_data_out_b_REG_field_type_0_sub_class_id; // @[XRam.scala 160:75]
  reg  io_data_out_b_REG_field_type_1_is_repeated; // @[XRam.scala 160:75]
  reg [4:0] io_data_out_b_REG_field_type_1_field_type; // @[XRam.scala 160:75]
  reg [15:0] io_data_out_b_REG_field_type_1_sub_class_id; // @[XRam.scala 160:75]
  reg  io_data_out_b_REG_field_type_2_is_repeated; // @[XRam.scala 160:75]
  reg [4:0] io_data_out_b_REG_field_type_2_field_type; // @[XRam.scala 160:75]
  reg [15:0] io_data_out_b_REG_field_type_2_sub_class_id; // @[XRam.scala 160:75]
  reg  io_data_out_b_REG_field_type_3_is_repeated; // @[XRam.scala 160:75]
  reg [4:0] io_data_out_b_REG_field_type_3_field_type; // @[XRam.scala 160:75]
  reg [15:0] io_data_out_b_REG_field_type_3_sub_class_id; // @[XRam.scala 160:75]
  reg  io_data_out_b_REG_field_type_4_is_repeated; // @[XRam.scala 160:75]
  reg [4:0] io_data_out_b_REG_field_type_4_field_type; // @[XRam.scala 160:75]
  reg [15:0] io_data_out_b_REG_field_type_4_sub_class_id; // @[XRam.scala 160:75]
  reg  io_data_out_b_REG_field_type_5_is_repeated; // @[XRam.scala 160:75]
  reg [4:0] io_data_out_b_REG_field_type_5_field_type; // @[XRam.scala 160:75]
  reg [15:0] io_data_out_b_REG_field_type_5_sub_class_id; // @[XRam.scala 160:75]
  reg  io_data_out_b_REG_field_type_6_is_repeated; // @[XRam.scala 160:75]
  reg [4:0] io_data_out_b_REG_field_type_6_field_type; // @[XRam.scala 160:75]
  reg [15:0] io_data_out_b_REG_field_type_6_sub_class_id; // @[XRam.scala 160:75]
  reg  io_data_out_b_REG_field_type_7_is_repeated; // @[XRam.scala 160:75]
  reg [4:0] io_data_out_b_REG_field_type_7_field_type; // @[XRam.scala 160:75]
  reg [15:0] io_data_out_b_REG_field_type_7_sub_class_id; // @[XRam.scala 160:75]
  reg  io_data_out_b_REG_field_type_8_is_repeated; // @[XRam.scala 160:75]
  reg [4:0] io_data_out_b_REG_field_type_8_field_type; // @[XRam.scala 160:75]
  reg [15:0] io_data_out_b_REG_field_type_8_sub_class_id; // @[XRam.scala 160:75]
  reg  io_data_out_b_REG_field_type_9_is_repeated; // @[XRam.scala 160:75]
  reg [4:0] io_data_out_b_REG_field_type_9_field_type; // @[XRam.scala 160:75]
  reg [15:0] io_data_out_b_REG_field_type_9_sub_class_id; // @[XRam.scala 160:75]
  reg  io_data_out_b_REG_field_type_10_is_repeated; // @[XRam.scala 160:75]
  reg [4:0] io_data_out_b_REG_field_type_10_field_type; // @[XRam.scala 160:75]
  reg [15:0] io_data_out_b_REG_field_type_10_sub_class_id; // @[XRam.scala 160:75]
  reg  io_data_out_b_REG_field_type_11_is_repeated; // @[XRam.scala 160:75]
  reg [4:0] io_data_out_b_REG_field_type_11_field_type; // @[XRam.scala 160:75]
  reg [15:0] io_data_out_b_REG_field_type_11_sub_class_id; // @[XRam.scala 160:75]
  reg  io_data_out_b_REG_field_type_12_is_repeated; // @[XRam.scala 160:75]
  reg [4:0] io_data_out_b_REG_field_type_12_field_type; // @[XRam.scala 160:75]
  reg [15:0] io_data_out_b_REG_field_type_12_sub_class_id; // @[XRam.scala 160:75]
  reg  io_data_out_b_REG_field_type_13_is_repeated; // @[XRam.scala 160:75]
  reg [4:0] io_data_out_b_REG_field_type_13_field_type; // @[XRam.scala 160:75]
  reg [15:0] io_data_out_b_REG_field_type_13_sub_class_id; // @[XRam.scala 160:75]
  reg  io_data_out_b_REG_field_type_14_is_repeated; // @[XRam.scala 160:75]
  reg [4:0] io_data_out_b_REG_field_type_14_field_type; // @[XRam.scala 160:75]
  reg [15:0] io_data_out_b_REG_field_type_14_sub_class_id; // @[XRam.scala 160:75]
  reg  io_data_out_b_REG_field_type_15_is_repeated; // @[XRam.scala 160:75]
  reg [4:0] io_data_out_b_REG_field_type_15_field_type; // @[XRam.scala 160:75]
  reg [15:0] io_data_out_b_REG_field_type_15_sub_class_id; // @[XRam.scala 160:75]
  reg  io_data_out_b_REG_field_type_16_is_repeated; // @[XRam.scala 160:75]
  reg [4:0] io_data_out_b_REG_field_type_16_field_type; // @[XRam.scala 160:75]
  reg [15:0] io_data_out_b_REG_field_type_16_sub_class_id; // @[XRam.scala 160:75]
  reg  io_data_out_b_REG_field_type_17_is_repeated; // @[XRam.scala 160:75]
  reg [4:0] io_data_out_b_REG_field_type_17_field_type; // @[XRam.scala 160:75]
  reg [15:0] io_data_out_b_REG_field_type_17_sub_class_id; // @[XRam.scala 160:75]
  reg  io_data_out_b_REG_field_type_18_is_repeated; // @[XRam.scala 160:75]
  reg [4:0] io_data_out_b_REG_field_type_18_field_type; // @[XRam.scala 160:75]
  reg [15:0] io_data_out_b_REG_field_type_18_sub_class_id; // @[XRam.scala 160:75]
  reg  io_data_out_b_REG_field_type_19_is_repeated; // @[XRam.scala 160:75]
  reg [4:0] io_data_out_b_REG_field_type_19_field_type; // @[XRam.scala 160:75]
  reg [15:0] io_data_out_b_REG_field_type_19_sub_class_id; // @[XRam.scala 160:75]
  reg  io_data_out_b_REG_field_type_20_is_repeated; // @[XRam.scala 160:75]
  reg [4:0] io_data_out_b_REG_field_type_20_field_type; // @[XRam.scala 160:75]
  reg [15:0] io_data_out_b_REG_field_type_20_sub_class_id; // @[XRam.scala 160:75]
  reg  io_data_out_b_REG_field_type_21_is_repeated; // @[XRam.scala 160:75]
  reg [4:0] io_data_out_b_REG_field_type_21_field_type; // @[XRam.scala 160:75]
  reg [15:0] io_data_out_b_REG_field_type_21_sub_class_id; // @[XRam.scala 160:75]
  reg  io_data_out_b_REG_field_type_22_is_repeated; // @[XRam.scala 160:75]
  reg [4:0] io_data_out_b_REG_field_type_22_field_type; // @[XRam.scala 160:75]
  reg [15:0] io_data_out_b_REG_field_type_22_sub_class_id; // @[XRam.scala 160:75]
  reg  io_data_out_b_REG_field_type_23_is_repeated; // @[XRam.scala 160:75]
  reg [4:0] io_data_out_b_REG_field_type_23_field_type; // @[XRam.scala 160:75]
  reg [15:0] io_data_out_b_REG_field_type_23_sub_class_id; // @[XRam.scala 160:75]
  reg  io_data_out_b_REG_field_type_24_is_repeated; // @[XRam.scala 160:75]
  reg [4:0] io_data_out_b_REG_field_type_24_field_type; // @[XRam.scala 160:75]
  reg [15:0] io_data_out_b_REG_field_type_24_sub_class_id; // @[XRam.scala 160:75]
  reg  io_data_out_b_REG_field_type_25_is_repeated; // @[XRam.scala 160:75]
  reg [4:0] io_data_out_b_REG_field_type_25_field_type; // @[XRam.scala 160:75]
  reg [15:0] io_data_out_b_REG_field_type_25_sub_class_id; // @[XRam.scala 160:75]
  reg  io_data_out_b_REG_field_type_26_is_repeated; // @[XRam.scala 160:75]
  reg [4:0] io_data_out_b_REG_field_type_26_field_type; // @[XRam.scala 160:75]
  reg [15:0] io_data_out_b_REG_field_type_26_sub_class_id; // @[XRam.scala 160:75]
  reg  io_data_out_b_REG_field_type_27_is_repeated; // @[XRam.scala 160:75]
  reg [4:0] io_data_out_b_REG_field_type_27_field_type; // @[XRam.scala 160:75]
  reg [15:0] io_data_out_b_REG_field_type_27_sub_class_id; // @[XRam.scala 160:75]
  reg  io_data_out_b_REG_field_type_28_is_repeated; // @[XRam.scala 160:75]
  reg [4:0] io_data_out_b_REG_field_type_28_field_type; // @[XRam.scala 160:75]
  reg [15:0] io_data_out_b_REG_field_type_28_sub_class_id; // @[XRam.scala 160:75]
  reg  io_data_out_b_REG_field_type_29_is_repeated; // @[XRam.scala 160:75]
  reg [4:0] io_data_out_b_REG_field_type_29_field_type; // @[XRam.scala 160:75]
  reg [15:0] io_data_out_b_REG_field_type_29_sub_class_id; // @[XRam.scala 160:75]
  reg  io_data_out_b_REG_field_type_30_is_repeated; // @[XRam.scala 160:75]
  reg [4:0] io_data_out_b_REG_field_type_30_field_type; // @[XRam.scala 160:75]
  reg [15:0] io_data_out_b_REG_field_type_30_sub_class_id; // @[XRam.scala 160:75]
  reg  io_data_out_b_REG_field_type_31_is_repeated; // @[XRam.scala 160:75]
  reg [4:0] io_data_out_b_REG_field_type_31_field_type; // @[XRam.scala 160:75]
  reg [15:0] io_data_out_b_REG_field_type_31_sub_class_id; // @[XRam.scala 160:75]
  reg  io_data_out_b_REG_field_type_32_is_repeated; // @[XRam.scala 160:75]
  reg [4:0] io_data_out_b_REG_field_type_32_field_type; // @[XRam.scala 160:75]
  reg [15:0] io_data_out_b_REG_field_type_32_sub_class_id; // @[XRam.scala 160:75]
  wire [45:0] ram_io_dina_lo_lo_lo_lo = {io_data_in_a_field_type_1_is_repeated,io_data_in_a_field_type_1_field_type,
    io_data_in_a_field_type_1_sub_class_id,io_data_in_a_field_type_1_is_host,io_data_in_a_field_type_0_is_repeated,
    io_data_in_a_field_type_0_field_type,io_data_in_a_field_type_0_sub_class_id,io_data_in_a_field_type_0_is_host}; // @[XRam.scala 184:106]
  wire [45:0] ram_io_dina_lo_lo_hi_lo = {io_data_in_a_field_type_5_is_repeated,io_data_in_a_field_type_5_field_type,
    io_data_in_a_field_type_5_sub_class_id,io_data_in_a_field_type_5_is_host,io_data_in_a_field_type_4_is_repeated,
    io_data_in_a_field_type_4_field_type,io_data_in_a_field_type_4_sub_class_id,io_data_in_a_field_type_4_is_host}; // @[XRam.scala 184:106]
  wire [92:0] ram_io_dina_lo_lo_hi = {io_data_in_a_field_type_8_is_host,io_data_in_a_field_type_7_is_repeated,
    io_data_in_a_field_type_7_field_type,io_data_in_a_field_type_7_sub_class_id,io_data_in_a_field_type_7_is_host,
    io_data_in_a_field_type_6_is_repeated,io_data_in_a_field_type_6_field_type,io_data_in_a_field_type_6_sub_class_id,
    io_data_in_a_field_type_6_is_host,ram_io_dina_lo_lo_hi_lo}; // @[XRam.scala 184:106]
  wire [184:0] ram_io_dina_lo_lo = {ram_io_dina_lo_lo_hi,io_data_in_a_field_type_3_is_repeated,
    io_data_in_a_field_type_3_field_type,io_data_in_a_field_type_3_sub_class_id,io_data_in_a_field_type_3_is_host,
    io_data_in_a_field_type_2_is_repeated,io_data_in_a_field_type_2_field_type,io_data_in_a_field_type_2_sub_class_id,
    io_data_in_a_field_type_2_is_host,ram_io_dina_lo_lo_lo_lo}; // @[XRam.scala 184:106]
  wire [45:0] ram_io_dina_lo_hi_lo_lo = {io_data_in_a_field_type_10_is_host,io_data_in_a_field_type_9_is_repeated,
    io_data_in_a_field_type_9_field_type,io_data_in_a_field_type_9_sub_class_id,io_data_in_a_field_type_9_is_host,
    io_data_in_a_field_type_8_is_repeated,io_data_in_a_field_type_8_field_type,io_data_in_a_field_type_8_sub_class_id}; // @[XRam.scala 184:106]
  wire [107:0] ram_io_dina_lo_hi_lo = {io_data_in_a_field_type_12_sub_class_id,io_data_in_a_field_type_12_is_host,
    io_data_in_a_field_type_11_is_repeated,io_data_in_a_field_type_11_field_type,io_data_in_a_field_type_11_sub_class_id
    ,io_data_in_a_field_type_11_is_host,io_data_in_a_field_type_10_is_repeated,io_data_in_a_field_type_10_field_type,
    io_data_in_a_field_type_10_sub_class_id,ram_io_dina_lo_hi_lo_lo}; // @[XRam.scala 184:106]
  wire [45:0] ram_io_dina_lo_hi_hi_lo = {io_data_in_a_field_type_14_sub_class_id,io_data_in_a_field_type_14_is_host,
    io_data_in_a_field_type_13_is_repeated,io_data_in_a_field_type_13_field_type,io_data_in_a_field_type_13_sub_class_id
    ,io_data_in_a_field_type_13_is_host,io_data_in_a_field_type_12_is_repeated,io_data_in_a_field_type_12_field_type}; // @[XRam.scala 184:106]
  wire [96:0] ram_io_dina_lo_hi_hi = {io_data_in_a_field_type_16_field_type,io_data_in_a_field_type_16_sub_class_id,
    io_data_in_a_field_type_16_is_host,io_data_in_a_field_type_15_is_repeated,io_data_in_a_field_type_15_field_type,
    io_data_in_a_field_type_15_sub_class_id,io_data_in_a_field_type_15_is_host,io_data_in_a_field_type_14_is_repeated,
    io_data_in_a_field_type_14_field_type,ram_io_dina_lo_hi_hi_lo}; // @[XRam.scala 184:106]
  wire [45:0] ram_io_dina_hi_lo_lo_lo = {io_data_in_a_field_type_18_field_type,io_data_in_a_field_type_18_sub_class_id,
    io_data_in_a_field_type_18_is_host,io_data_in_a_field_type_17_is_repeated,io_data_in_a_field_type_17_field_type,
    io_data_in_a_field_type_17_sub_class_id,io_data_in_a_field_type_17_is_host,io_data_in_a_field_type_16_is_repeated}; // @[XRam.scala 184:106]
  wire [45:0] ram_io_dina_hi_lo_hi_lo = {io_data_in_a_field_type_22_field_type,io_data_in_a_field_type_22_sub_class_id,
    io_data_in_a_field_type_22_is_host,io_data_in_a_field_type_21_is_repeated,io_data_in_a_field_type_21_field_type,
    io_data_in_a_field_type_21_sub_class_id,io_data_in_a_field_type_21_is_host,io_data_in_a_field_type_20_is_repeated}; // @[XRam.scala 184:106]
  wire [92:0] ram_io_dina_hi_lo_hi = {io_data_in_a_field_type_24_is_repeated,io_data_in_a_field_type_24_field_type,
    io_data_in_a_field_type_24_sub_class_id,io_data_in_a_field_type_24_is_host,io_data_in_a_field_type_23_is_repeated,
    io_data_in_a_field_type_23_field_type,io_data_in_a_field_type_23_sub_class_id,io_data_in_a_field_type_23_is_host,
    io_data_in_a_field_type_22_is_repeated,ram_io_dina_hi_lo_hi_lo}; // @[XRam.scala 184:106]
  wire [184:0] ram_io_dina_hi_lo = {ram_io_dina_hi_lo_hi,io_data_in_a_field_type_20_field_type,
    io_data_in_a_field_type_20_sub_class_id,io_data_in_a_field_type_20_is_host,io_data_in_a_field_type_19_is_repeated,
    io_data_in_a_field_type_19_field_type,io_data_in_a_field_type_19_sub_class_id,io_data_in_a_field_type_19_is_host,
    io_data_in_a_field_type_18_is_repeated,ram_io_dina_hi_lo_lo_lo}; // @[XRam.scala 184:106]
  wire [45:0] ram_io_dina_hi_hi_lo_lo = {io_data_in_a_field_type_26_is_repeated,io_data_in_a_field_type_26_field_type,
    io_data_in_a_field_type_26_sub_class_id,io_data_in_a_field_type_26_is_host,io_data_in_a_field_type_25_is_repeated,
    io_data_in_a_field_type_25_field_type,io_data_in_a_field_type_25_sub_class_id,io_data_in_a_field_type_25_is_host}; // @[XRam.scala 184:106]
  wire [92:0] ram_io_dina_hi_hi_lo = {io_data_in_a_field_type_29_is_host,io_data_in_a_field_type_28_is_repeated,
    io_data_in_a_field_type_28_field_type,io_data_in_a_field_type_28_sub_class_id,io_data_in_a_field_type_28_is_host,
    io_data_in_a_field_type_27_is_repeated,io_data_in_a_field_type_27_field_type,io_data_in_a_field_type_27_sub_class_id
    ,io_data_in_a_field_type_27_is_host,ram_io_dina_hi_hi_lo_lo}; // @[XRam.scala 184:106]
  wire [45:0] ram_io_dina_hi_hi_hi_lo = {io_data_in_a_field_type_31_is_host,io_data_in_a_field_type_30_is_repeated,
    io_data_in_a_field_type_30_field_type,io_data_in_a_field_type_30_sub_class_id,io_data_in_a_field_type_30_is_host,
    io_data_in_a_field_type_29_is_repeated,io_data_in_a_field_type_29_field_type,io_data_in_a_field_type_29_sub_class_id
    }; // @[XRam.scala 184:106]
  wire [114:0] ram_io_dina_hi_hi_hi = {io_data_in_a_class_length,io_data_in_a_max_field_num,
    io_data_in_a_field_type_32_is_repeated,io_data_in_a_field_type_32_field_type,io_data_in_a_field_type_32_sub_class_id
    ,io_data_in_a_field_type_32_is_host,io_data_in_a_field_type_31_is_repeated,io_data_in_a_field_type_31_field_type,
    io_data_in_a_field_type_31_sub_class_id,ram_io_dina_hi_hi_hi_lo}; // @[XRam.scala 184:106]
  wire [782:0] _ram_io_dina_T_1 = {ram_io_dina_hi_hi_hi,ram_io_dina_hi_hi_lo,ram_io_dina_hi_lo,ram_io_dina_lo_hi_hi,
    ram_io_dina_lo_hi_lo,ram_io_dina_lo_lo}; // @[XRam.scala 184:106]
  wire [782:0] _ram_io_dina_T_2 = usr_rst_delay ? 783'h0 : _ram_io_dina_T_1; // @[XRam.scala 184:63]
  xpm_memory_tdpram
    #(.USE_EMBEDDED_CONSTRAINT(0), .CLOCKING_MODE("common_clock"), .WRITE_DATA_WIDTH_B(784), .READ_LATENCY_B(1), .ADDR_WIDTH_A(10), .READ_DATA_WIDTH_A(784), .RST_MODE_B("SYNC"), .WAKEUP_TIME("disable_sleep"), .MEMORY_INIT_FILE("none"), .READ_LATENCY_A(1), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_A(784), .AUTO_SLEEP_TIME(0), .WRITE_MODE_A("no_change"), .MEMORY_PRIMITIVE("auto"), .USE_MEM_INIT(1), .MEMORY_INIT_PARAM(""), .SIM_ASSERT_CHK(0), .ECC_MODE("no_ecc"), .READ_RESET_VALUE_A("0"), .BYTE_WRITE_WIDTH_A(8), .MEMORY_OPTIMIZATION("true"), .MESSAGE_CONTROL(0), .WRITE_MODE_B("no_change"), .READ_DATA_WIDTH_B(784), .ADDR_WIDTH_B(10), .CASCADE_HEIGHT(0), .READ_RESET_VALUE_B("0"), .BYTE_WRITE_WIDTH_B(8), .MEMORY_SIZE(802816))
    ram ( // @[XRam.scala 136:33]
    .douta(ram_douta),
    .doutb(ram_doutb),
    .addra(ram_addra),
    .addrb(ram_addrb),
    .clka(ram_clka),
    .clkb(ram_clkb),
    .dina(ram_dina),
    .dinb(ram_dinb),
    .ena(ram_ena),
    .enb(ram_enb),
    .injectdbiterra(ram_injectdbiterra),
    .injectdbiterrb(ram_injectdbiterrb),
    .injectsbiterra(ram_injectsbiterra),
    .injectsbiterrb(ram_injectsbiterrb),
    .regcea(ram_regcea),
    .regceb(ram_regceb),
    .rsta(ram_rsta),
    .rstb(ram_rstb),
    .sleep(ram_sleep),
    .wea(ram_wea),
    .web(ram_web)
  );
  assign io_data_out_b_max_field_num = REG == REG_1 & REG_2 ? io_data_out_b_REG_max_field_num : ram_doutb[766:759]; // @[XRam.scala 159:102 XRam.scala 160:65 XRam.scala 162:65]
  assign io_data_out_b_field_type_0_is_repeated = REG == REG_1 & REG_2 ? io_data_out_b_REG_field_type_0_is_repeated :
    ram_doutb[22]; // @[XRam.scala 159:102 XRam.scala 160:65 XRam.scala 162:65]
  assign io_data_out_b_field_type_0_field_type = REG == REG_1 & REG_2 ? io_data_out_b_REG_field_type_0_field_type :
    ram_doutb[21:17]; // @[XRam.scala 159:102 XRam.scala 160:65 XRam.scala 162:65]
  assign io_data_out_b_field_type_0_sub_class_id = REG == REG_1 & REG_2 ? io_data_out_b_REG_field_type_0_sub_class_id :
    ram_doutb[16:1]; // @[XRam.scala 159:102 XRam.scala 160:65 XRam.scala 162:65]
  assign io_data_out_b_field_type_1_is_repeated = REG == REG_1 & REG_2 ? io_data_out_b_REG_field_type_1_is_repeated :
    ram_doutb[45]; // @[XRam.scala 159:102 XRam.scala 160:65 XRam.scala 162:65]
  assign io_data_out_b_field_type_1_field_type = REG == REG_1 & REG_2 ? io_data_out_b_REG_field_type_1_field_type :
    ram_doutb[44:40]; // @[XRam.scala 159:102 XRam.scala 160:65 XRam.scala 162:65]
  assign io_data_out_b_field_type_1_sub_class_id = REG == REG_1 & REG_2 ? io_data_out_b_REG_field_type_1_sub_class_id :
    ram_doutb[39:24]; // @[XRam.scala 159:102 XRam.scala 160:65 XRam.scala 162:65]
  assign io_data_out_b_field_type_2_is_repeated = REG == REG_1 & REG_2 ? io_data_out_b_REG_field_type_2_is_repeated :
    ram_doutb[68]; // @[XRam.scala 159:102 XRam.scala 160:65 XRam.scala 162:65]
  assign io_data_out_b_field_type_2_field_type = REG == REG_1 & REG_2 ? io_data_out_b_REG_field_type_2_field_type :
    ram_doutb[67:63]; // @[XRam.scala 159:102 XRam.scala 160:65 XRam.scala 162:65]
  assign io_data_out_b_field_type_2_sub_class_id = REG == REG_1 & REG_2 ? io_data_out_b_REG_field_type_2_sub_class_id :
    ram_doutb[62:47]; // @[XRam.scala 159:102 XRam.scala 160:65 XRam.scala 162:65]
  assign io_data_out_b_field_type_3_is_repeated = REG == REG_1 & REG_2 ? io_data_out_b_REG_field_type_3_is_repeated :
    ram_doutb[91]; // @[XRam.scala 159:102 XRam.scala 160:65 XRam.scala 162:65]
  assign io_data_out_b_field_type_3_field_type = REG == REG_1 & REG_2 ? io_data_out_b_REG_field_type_3_field_type :
    ram_doutb[90:86]; // @[XRam.scala 159:102 XRam.scala 160:65 XRam.scala 162:65]
  assign io_data_out_b_field_type_3_sub_class_id = REG == REG_1 & REG_2 ? io_data_out_b_REG_field_type_3_sub_class_id :
    ram_doutb[85:70]; // @[XRam.scala 159:102 XRam.scala 160:65 XRam.scala 162:65]
  assign io_data_out_b_field_type_4_is_repeated = REG == REG_1 & REG_2 ? io_data_out_b_REG_field_type_4_is_repeated :
    ram_doutb[114]; // @[XRam.scala 159:102 XRam.scala 160:65 XRam.scala 162:65]
  assign io_data_out_b_field_type_4_field_type = REG == REG_1 & REG_2 ? io_data_out_b_REG_field_type_4_field_type :
    ram_doutb[113:109]; // @[XRam.scala 159:102 XRam.scala 160:65 XRam.scala 162:65]
  assign io_data_out_b_field_type_4_sub_class_id = REG == REG_1 & REG_2 ? io_data_out_b_REG_field_type_4_sub_class_id :
    ram_doutb[108:93]; // @[XRam.scala 159:102 XRam.scala 160:65 XRam.scala 162:65]
  assign io_data_out_b_field_type_5_is_repeated = REG == REG_1 & REG_2 ? io_data_out_b_REG_field_type_5_is_repeated :
    ram_doutb[137]; // @[XRam.scala 159:102 XRam.scala 160:65 XRam.scala 162:65]
  assign io_data_out_b_field_type_5_field_type = REG == REG_1 & REG_2 ? io_data_out_b_REG_field_type_5_field_type :
    ram_doutb[136:132]; // @[XRam.scala 159:102 XRam.scala 160:65 XRam.scala 162:65]
  assign io_data_out_b_field_type_5_sub_class_id = REG == REG_1 & REG_2 ? io_data_out_b_REG_field_type_5_sub_class_id :
    ram_doutb[131:116]; // @[XRam.scala 159:102 XRam.scala 160:65 XRam.scala 162:65]
  assign io_data_out_b_field_type_6_is_repeated = REG == REG_1 & REG_2 ? io_data_out_b_REG_field_type_6_is_repeated :
    ram_doutb[160]; // @[XRam.scala 159:102 XRam.scala 160:65 XRam.scala 162:65]
  assign io_data_out_b_field_type_6_field_type = REG == REG_1 & REG_2 ? io_data_out_b_REG_field_type_6_field_type :
    ram_doutb[159:155]; // @[XRam.scala 159:102 XRam.scala 160:65 XRam.scala 162:65]
  assign io_data_out_b_field_type_6_sub_class_id = REG == REG_1 & REG_2 ? io_data_out_b_REG_field_type_6_sub_class_id :
    ram_doutb[154:139]; // @[XRam.scala 159:102 XRam.scala 160:65 XRam.scala 162:65]
  assign io_data_out_b_field_type_7_is_repeated = REG == REG_1 & REG_2 ? io_data_out_b_REG_field_type_7_is_repeated :
    ram_doutb[183]; // @[XRam.scala 159:102 XRam.scala 160:65 XRam.scala 162:65]
  assign io_data_out_b_field_type_7_field_type = REG == REG_1 & REG_2 ? io_data_out_b_REG_field_type_7_field_type :
    ram_doutb[182:178]; // @[XRam.scala 159:102 XRam.scala 160:65 XRam.scala 162:65]
  assign io_data_out_b_field_type_7_sub_class_id = REG == REG_1 & REG_2 ? io_data_out_b_REG_field_type_7_sub_class_id :
    ram_doutb[177:162]; // @[XRam.scala 159:102 XRam.scala 160:65 XRam.scala 162:65]
  assign io_data_out_b_field_type_8_is_repeated = REG == REG_1 & REG_2 ? io_data_out_b_REG_field_type_8_is_repeated :
    ram_doutb[206]; // @[XRam.scala 159:102 XRam.scala 160:65 XRam.scala 162:65]
  assign io_data_out_b_field_type_8_field_type = REG == REG_1 & REG_2 ? io_data_out_b_REG_field_type_8_field_type :
    ram_doutb[205:201]; // @[XRam.scala 159:102 XRam.scala 160:65 XRam.scala 162:65]
  assign io_data_out_b_field_type_8_sub_class_id = REG == REG_1 & REG_2 ? io_data_out_b_REG_field_type_8_sub_class_id :
    ram_doutb[200:185]; // @[XRam.scala 159:102 XRam.scala 160:65 XRam.scala 162:65]
  assign io_data_out_b_field_type_9_is_repeated = REG == REG_1 & REG_2 ? io_data_out_b_REG_field_type_9_is_repeated :
    ram_doutb[229]; // @[XRam.scala 159:102 XRam.scala 160:65 XRam.scala 162:65]
  assign io_data_out_b_field_type_9_field_type = REG == REG_1 & REG_2 ? io_data_out_b_REG_field_type_9_field_type :
    ram_doutb[228:224]; // @[XRam.scala 159:102 XRam.scala 160:65 XRam.scala 162:65]
  assign io_data_out_b_field_type_9_sub_class_id = REG == REG_1 & REG_2 ? io_data_out_b_REG_field_type_9_sub_class_id :
    ram_doutb[223:208]; // @[XRam.scala 159:102 XRam.scala 160:65 XRam.scala 162:65]
  assign io_data_out_b_field_type_10_is_repeated = REG == REG_1 & REG_2 ? io_data_out_b_REG_field_type_10_is_repeated :
    ram_doutb[252]; // @[XRam.scala 159:102 XRam.scala 160:65 XRam.scala 162:65]
  assign io_data_out_b_field_type_10_field_type = REG == REG_1 & REG_2 ? io_data_out_b_REG_field_type_10_field_type :
    ram_doutb[251:247]; // @[XRam.scala 159:102 XRam.scala 160:65 XRam.scala 162:65]
  assign io_data_out_b_field_type_10_sub_class_id = REG == REG_1 & REG_2 ? io_data_out_b_REG_field_type_10_sub_class_id
     : ram_doutb[246:231]; // @[XRam.scala 159:102 XRam.scala 160:65 XRam.scala 162:65]
  assign io_data_out_b_field_type_11_is_repeated = REG == REG_1 & REG_2 ? io_data_out_b_REG_field_type_11_is_repeated :
    ram_doutb[275]; // @[XRam.scala 159:102 XRam.scala 160:65 XRam.scala 162:65]
  assign io_data_out_b_field_type_11_field_type = REG == REG_1 & REG_2 ? io_data_out_b_REG_field_type_11_field_type :
    ram_doutb[274:270]; // @[XRam.scala 159:102 XRam.scala 160:65 XRam.scala 162:65]
  assign io_data_out_b_field_type_11_sub_class_id = REG == REG_1 & REG_2 ? io_data_out_b_REG_field_type_11_sub_class_id
     : ram_doutb[269:254]; // @[XRam.scala 159:102 XRam.scala 160:65 XRam.scala 162:65]
  assign io_data_out_b_field_type_12_is_repeated = REG == REG_1 & REG_2 ? io_data_out_b_REG_field_type_12_is_repeated :
    ram_doutb[298]; // @[XRam.scala 159:102 XRam.scala 160:65 XRam.scala 162:65]
  assign io_data_out_b_field_type_12_field_type = REG == REG_1 & REG_2 ? io_data_out_b_REG_field_type_12_field_type :
    ram_doutb[297:293]; // @[XRam.scala 159:102 XRam.scala 160:65 XRam.scala 162:65]
  assign io_data_out_b_field_type_12_sub_class_id = REG == REG_1 & REG_2 ? io_data_out_b_REG_field_type_12_sub_class_id
     : ram_doutb[292:277]; // @[XRam.scala 159:102 XRam.scala 160:65 XRam.scala 162:65]
  assign io_data_out_b_field_type_13_is_repeated = REG == REG_1 & REG_2 ? io_data_out_b_REG_field_type_13_is_repeated :
    ram_doutb[321]; // @[XRam.scala 159:102 XRam.scala 160:65 XRam.scala 162:65]
  assign io_data_out_b_field_type_13_field_type = REG == REG_1 & REG_2 ? io_data_out_b_REG_field_type_13_field_type :
    ram_doutb[320:316]; // @[XRam.scala 159:102 XRam.scala 160:65 XRam.scala 162:65]
  assign io_data_out_b_field_type_13_sub_class_id = REG == REG_1 & REG_2 ? io_data_out_b_REG_field_type_13_sub_class_id
     : ram_doutb[315:300]; // @[XRam.scala 159:102 XRam.scala 160:65 XRam.scala 162:65]
  assign io_data_out_b_field_type_14_is_repeated = REG == REG_1 & REG_2 ? io_data_out_b_REG_field_type_14_is_repeated :
    ram_doutb[344]; // @[XRam.scala 159:102 XRam.scala 160:65 XRam.scala 162:65]
  assign io_data_out_b_field_type_14_field_type = REG == REG_1 & REG_2 ? io_data_out_b_REG_field_type_14_field_type :
    ram_doutb[343:339]; // @[XRam.scala 159:102 XRam.scala 160:65 XRam.scala 162:65]
  assign io_data_out_b_field_type_14_sub_class_id = REG == REG_1 & REG_2 ? io_data_out_b_REG_field_type_14_sub_class_id
     : ram_doutb[338:323]; // @[XRam.scala 159:102 XRam.scala 160:65 XRam.scala 162:65]
  assign io_data_out_b_field_type_15_is_repeated = REG == REG_1 & REG_2 ? io_data_out_b_REG_field_type_15_is_repeated :
    ram_doutb[367]; // @[XRam.scala 159:102 XRam.scala 160:65 XRam.scala 162:65]
  assign io_data_out_b_field_type_15_field_type = REG == REG_1 & REG_2 ? io_data_out_b_REG_field_type_15_field_type :
    ram_doutb[366:362]; // @[XRam.scala 159:102 XRam.scala 160:65 XRam.scala 162:65]
  assign io_data_out_b_field_type_15_sub_class_id = REG == REG_1 & REG_2 ? io_data_out_b_REG_field_type_15_sub_class_id
     : ram_doutb[361:346]; // @[XRam.scala 159:102 XRam.scala 160:65 XRam.scala 162:65]
  assign io_data_out_b_field_type_16_is_repeated = REG == REG_1 & REG_2 ? io_data_out_b_REG_field_type_16_is_repeated :
    ram_doutb[390]; // @[XRam.scala 159:102 XRam.scala 160:65 XRam.scala 162:65]
  assign io_data_out_b_field_type_16_field_type = REG == REG_1 & REG_2 ? io_data_out_b_REG_field_type_16_field_type :
    ram_doutb[389:385]; // @[XRam.scala 159:102 XRam.scala 160:65 XRam.scala 162:65]
  assign io_data_out_b_field_type_16_sub_class_id = REG == REG_1 & REG_2 ? io_data_out_b_REG_field_type_16_sub_class_id
     : ram_doutb[384:369]; // @[XRam.scala 159:102 XRam.scala 160:65 XRam.scala 162:65]
  assign io_data_out_b_field_type_17_is_repeated = REG == REG_1 & REG_2 ? io_data_out_b_REG_field_type_17_is_repeated :
    ram_doutb[413]; // @[XRam.scala 159:102 XRam.scala 160:65 XRam.scala 162:65]
  assign io_data_out_b_field_type_17_field_type = REG == REG_1 & REG_2 ? io_data_out_b_REG_field_type_17_field_type :
    ram_doutb[412:408]; // @[XRam.scala 159:102 XRam.scala 160:65 XRam.scala 162:65]
  assign io_data_out_b_field_type_17_sub_class_id = REG == REG_1 & REG_2 ? io_data_out_b_REG_field_type_17_sub_class_id
     : ram_doutb[407:392]; // @[XRam.scala 159:102 XRam.scala 160:65 XRam.scala 162:65]
  assign io_data_out_b_field_type_18_is_repeated = REG == REG_1 & REG_2 ? io_data_out_b_REG_field_type_18_is_repeated :
    ram_doutb[436]; // @[XRam.scala 159:102 XRam.scala 160:65 XRam.scala 162:65]
  assign io_data_out_b_field_type_18_field_type = REG == REG_1 & REG_2 ? io_data_out_b_REG_field_type_18_field_type :
    ram_doutb[435:431]; // @[XRam.scala 159:102 XRam.scala 160:65 XRam.scala 162:65]
  assign io_data_out_b_field_type_18_sub_class_id = REG == REG_1 & REG_2 ? io_data_out_b_REG_field_type_18_sub_class_id
     : ram_doutb[430:415]; // @[XRam.scala 159:102 XRam.scala 160:65 XRam.scala 162:65]
  assign io_data_out_b_field_type_19_is_repeated = REG == REG_1 & REG_2 ? io_data_out_b_REG_field_type_19_is_repeated :
    ram_doutb[459]; // @[XRam.scala 159:102 XRam.scala 160:65 XRam.scala 162:65]
  assign io_data_out_b_field_type_19_field_type = REG == REG_1 & REG_2 ? io_data_out_b_REG_field_type_19_field_type :
    ram_doutb[458:454]; // @[XRam.scala 159:102 XRam.scala 160:65 XRam.scala 162:65]
  assign io_data_out_b_field_type_19_sub_class_id = REG == REG_1 & REG_2 ? io_data_out_b_REG_field_type_19_sub_class_id
     : ram_doutb[453:438]; // @[XRam.scala 159:102 XRam.scala 160:65 XRam.scala 162:65]
  assign io_data_out_b_field_type_20_is_repeated = REG == REG_1 & REG_2 ? io_data_out_b_REG_field_type_20_is_repeated :
    ram_doutb[482]; // @[XRam.scala 159:102 XRam.scala 160:65 XRam.scala 162:65]
  assign io_data_out_b_field_type_20_field_type = REG == REG_1 & REG_2 ? io_data_out_b_REG_field_type_20_field_type :
    ram_doutb[481:477]; // @[XRam.scala 159:102 XRam.scala 160:65 XRam.scala 162:65]
  assign io_data_out_b_field_type_20_sub_class_id = REG == REG_1 & REG_2 ? io_data_out_b_REG_field_type_20_sub_class_id
     : ram_doutb[476:461]; // @[XRam.scala 159:102 XRam.scala 160:65 XRam.scala 162:65]
  assign io_data_out_b_field_type_21_is_repeated = REG == REG_1 & REG_2 ? io_data_out_b_REG_field_type_21_is_repeated :
    ram_doutb[505]; // @[XRam.scala 159:102 XRam.scala 160:65 XRam.scala 162:65]
  assign io_data_out_b_field_type_21_field_type = REG == REG_1 & REG_2 ? io_data_out_b_REG_field_type_21_field_type :
    ram_doutb[504:500]; // @[XRam.scala 159:102 XRam.scala 160:65 XRam.scala 162:65]
  assign io_data_out_b_field_type_21_sub_class_id = REG == REG_1 & REG_2 ? io_data_out_b_REG_field_type_21_sub_class_id
     : ram_doutb[499:484]; // @[XRam.scala 159:102 XRam.scala 160:65 XRam.scala 162:65]
  assign io_data_out_b_field_type_22_is_repeated = REG == REG_1 & REG_2 ? io_data_out_b_REG_field_type_22_is_repeated :
    ram_doutb[528]; // @[XRam.scala 159:102 XRam.scala 160:65 XRam.scala 162:65]
  assign io_data_out_b_field_type_22_field_type = REG == REG_1 & REG_2 ? io_data_out_b_REG_field_type_22_field_type :
    ram_doutb[527:523]; // @[XRam.scala 159:102 XRam.scala 160:65 XRam.scala 162:65]
  assign io_data_out_b_field_type_22_sub_class_id = REG == REG_1 & REG_2 ? io_data_out_b_REG_field_type_22_sub_class_id
     : ram_doutb[522:507]; // @[XRam.scala 159:102 XRam.scala 160:65 XRam.scala 162:65]
  assign io_data_out_b_field_type_23_is_repeated = REG == REG_1 & REG_2 ? io_data_out_b_REG_field_type_23_is_repeated :
    ram_doutb[551]; // @[XRam.scala 159:102 XRam.scala 160:65 XRam.scala 162:65]
  assign io_data_out_b_field_type_23_field_type = REG == REG_1 & REG_2 ? io_data_out_b_REG_field_type_23_field_type :
    ram_doutb[550:546]; // @[XRam.scala 159:102 XRam.scala 160:65 XRam.scala 162:65]
  assign io_data_out_b_field_type_23_sub_class_id = REG == REG_1 & REG_2 ? io_data_out_b_REG_field_type_23_sub_class_id
     : ram_doutb[545:530]; // @[XRam.scala 159:102 XRam.scala 160:65 XRam.scala 162:65]
  assign io_data_out_b_field_type_24_is_repeated = REG == REG_1 & REG_2 ? io_data_out_b_REG_field_type_24_is_repeated :
    ram_doutb[574]; // @[XRam.scala 159:102 XRam.scala 160:65 XRam.scala 162:65]
  assign io_data_out_b_field_type_24_field_type = REG == REG_1 & REG_2 ? io_data_out_b_REG_field_type_24_field_type :
    ram_doutb[573:569]; // @[XRam.scala 159:102 XRam.scala 160:65 XRam.scala 162:65]
  assign io_data_out_b_field_type_24_sub_class_id = REG == REG_1 & REG_2 ? io_data_out_b_REG_field_type_24_sub_class_id
     : ram_doutb[568:553]; // @[XRam.scala 159:102 XRam.scala 160:65 XRam.scala 162:65]
  assign io_data_out_b_field_type_25_is_repeated = REG == REG_1 & REG_2 ? io_data_out_b_REG_field_type_25_is_repeated :
    ram_doutb[597]; // @[XRam.scala 159:102 XRam.scala 160:65 XRam.scala 162:65]
  assign io_data_out_b_field_type_25_field_type = REG == REG_1 & REG_2 ? io_data_out_b_REG_field_type_25_field_type :
    ram_doutb[596:592]; // @[XRam.scala 159:102 XRam.scala 160:65 XRam.scala 162:65]
  assign io_data_out_b_field_type_25_sub_class_id = REG == REG_1 & REG_2 ? io_data_out_b_REG_field_type_25_sub_class_id
     : ram_doutb[591:576]; // @[XRam.scala 159:102 XRam.scala 160:65 XRam.scala 162:65]
  assign io_data_out_b_field_type_26_is_repeated = REG == REG_1 & REG_2 ? io_data_out_b_REG_field_type_26_is_repeated :
    ram_doutb[620]; // @[XRam.scala 159:102 XRam.scala 160:65 XRam.scala 162:65]
  assign io_data_out_b_field_type_26_field_type = REG == REG_1 & REG_2 ? io_data_out_b_REG_field_type_26_field_type :
    ram_doutb[619:615]; // @[XRam.scala 159:102 XRam.scala 160:65 XRam.scala 162:65]
  assign io_data_out_b_field_type_26_sub_class_id = REG == REG_1 & REG_2 ? io_data_out_b_REG_field_type_26_sub_class_id
     : ram_doutb[614:599]; // @[XRam.scala 159:102 XRam.scala 160:65 XRam.scala 162:65]
  assign io_data_out_b_field_type_27_is_repeated = REG == REG_1 & REG_2 ? io_data_out_b_REG_field_type_27_is_repeated :
    ram_doutb[643]; // @[XRam.scala 159:102 XRam.scala 160:65 XRam.scala 162:65]
  assign io_data_out_b_field_type_27_field_type = REG == REG_1 & REG_2 ? io_data_out_b_REG_field_type_27_field_type :
    ram_doutb[642:638]; // @[XRam.scala 159:102 XRam.scala 160:65 XRam.scala 162:65]
  assign io_data_out_b_field_type_27_sub_class_id = REG == REG_1 & REG_2 ? io_data_out_b_REG_field_type_27_sub_class_id
     : ram_doutb[637:622]; // @[XRam.scala 159:102 XRam.scala 160:65 XRam.scala 162:65]
  assign io_data_out_b_field_type_28_is_repeated = REG == REG_1 & REG_2 ? io_data_out_b_REG_field_type_28_is_repeated :
    ram_doutb[666]; // @[XRam.scala 159:102 XRam.scala 160:65 XRam.scala 162:65]
  assign io_data_out_b_field_type_28_field_type = REG == REG_1 & REG_2 ? io_data_out_b_REG_field_type_28_field_type :
    ram_doutb[665:661]; // @[XRam.scala 159:102 XRam.scala 160:65 XRam.scala 162:65]
  assign io_data_out_b_field_type_28_sub_class_id = REG == REG_1 & REG_2 ? io_data_out_b_REG_field_type_28_sub_class_id
     : ram_doutb[660:645]; // @[XRam.scala 159:102 XRam.scala 160:65 XRam.scala 162:65]
  assign io_data_out_b_field_type_29_is_repeated = REG == REG_1 & REG_2 ? io_data_out_b_REG_field_type_29_is_repeated :
    ram_doutb[689]; // @[XRam.scala 159:102 XRam.scala 160:65 XRam.scala 162:65]
  assign io_data_out_b_field_type_29_field_type = REG == REG_1 & REG_2 ? io_data_out_b_REG_field_type_29_field_type :
    ram_doutb[688:684]; // @[XRam.scala 159:102 XRam.scala 160:65 XRam.scala 162:65]
  assign io_data_out_b_field_type_29_sub_class_id = REG == REG_1 & REG_2 ? io_data_out_b_REG_field_type_29_sub_class_id
     : ram_doutb[683:668]; // @[XRam.scala 159:102 XRam.scala 160:65 XRam.scala 162:65]
  assign io_data_out_b_field_type_30_is_repeated = REG == REG_1 & REG_2 ? io_data_out_b_REG_field_type_30_is_repeated :
    ram_doutb[712]; // @[XRam.scala 159:102 XRam.scala 160:65 XRam.scala 162:65]
  assign io_data_out_b_field_type_30_field_type = REG == REG_1 & REG_2 ? io_data_out_b_REG_field_type_30_field_type :
    ram_doutb[711:707]; // @[XRam.scala 159:102 XRam.scala 160:65 XRam.scala 162:65]
  assign io_data_out_b_field_type_30_sub_class_id = REG == REG_1 & REG_2 ? io_data_out_b_REG_field_type_30_sub_class_id
     : ram_doutb[706:691]; // @[XRam.scala 159:102 XRam.scala 160:65 XRam.scala 162:65]
  assign io_data_out_b_field_type_31_is_repeated = REG == REG_1 & REG_2 ? io_data_out_b_REG_field_type_31_is_repeated :
    ram_doutb[735]; // @[XRam.scala 159:102 XRam.scala 160:65 XRam.scala 162:65]
  assign io_data_out_b_field_type_31_field_type = REG == REG_1 & REG_2 ? io_data_out_b_REG_field_type_31_field_type :
    ram_doutb[734:730]; // @[XRam.scala 159:102 XRam.scala 160:65 XRam.scala 162:65]
  assign io_data_out_b_field_type_31_sub_class_id = REG == REG_1 & REG_2 ? io_data_out_b_REG_field_type_31_sub_class_id
     : ram_doutb[729:714]; // @[XRam.scala 159:102 XRam.scala 160:65 XRam.scala 162:65]
  assign io_data_out_b_field_type_32_is_repeated = REG == REG_1 & REG_2 ? io_data_out_b_REG_field_type_32_is_repeated :
    ram_doutb[758]; // @[XRam.scala 159:102 XRam.scala 160:65 XRam.scala 162:65]
  assign io_data_out_b_field_type_32_field_type = REG == REG_1 & REG_2 ? io_data_out_b_REG_field_type_32_field_type :
    ram_doutb[757:753]; // @[XRam.scala 159:102 XRam.scala 160:65 XRam.scala 162:65]
  assign io_data_out_b_field_type_32_sub_class_id = REG == REG_1 & REG_2 ? io_data_out_b_REG_field_type_32_sub_class_id
     : ram_doutb[752:737]; // @[XRam.scala 159:102 XRam.scala 160:65 XRam.scala 162:65]
  assign ram_addra = usr_rst_delay ? reset_addr : io_addr_a; // @[XRam.scala 178:55]
  assign ram_addrb = io_addr_b; // @[XRam.scala 179:49]
  assign ram_clka = clock; // @[XRam.scala 181:57]
  assign ram_clkb = clock; // @[XRam.scala 182:57]
  assign ram_dina = {{1'd0}, _ram_io_dina_T_2}; // @[XRam.scala 184:63]
  assign ram_dinb = 784'h0; // @[XRam.scala 185:57]
  assign ram_ena = 1'h1; // @[XRam.scala 187:57]
  assign ram_enb = 1'h1; // @[XRam.scala 188:57]
  assign ram_injectdbiterra = 1'h0; // @[XRam.scala 190:41]
  assign ram_injectdbiterrb = 1'h0; // @[XRam.scala 191:41]
  assign ram_injectsbiterra = 1'h0; // @[XRam.scala 193:41]
  assign ram_injectsbiterrb = 1'h0; // @[XRam.scala 194:41]
  assign ram_regcea = 1'h1; // @[XRam.scala 196:49]
  assign ram_regceb = 1'h1; // @[XRam.scala 197:49]
  assign ram_rsta = 1'h0; // @[XRam.scala 199:57]
  assign ram_rstb = 1'h0; // @[XRam.scala 200:57]
  assign ram_sleep = 1'h0; // @[XRam.scala 202:49]
  assign ram_wea = usr_rst_delay ? 98'h3ffffffffffffffffffffffff : wr_en_a; // @[XRam.scala 206:63]
  assign ram_web = 98'h0; // @[XRam.scala 208:57]
  always @(posedge clock) begin
    usr_rst_delay_r <= reset; // @[Reg.scala 16:19 Reg.scala 16:23 Reg.scala 15:16]
    usr_rst_delay_r_1 <= usr_rst_delay_r; // @[Reg.scala 16:19 Reg.scala 16:23 Reg.scala 15:16]
    usr_rst_delay_r_2 <= usr_rst_delay_r_1; // @[Reg.scala 16:19 Reg.scala 16:23 Reg.scala 15:16]
    usr_rst_delay <= usr_rst_delay_r_2; // @[Reg.scala 16:19 Reg.scala 16:23 Reg.scala 15:16]
    if (usr_rst_delay) begin // @[XRam.scala 143:45]
      reset_addr <= _reset_addr_T_1; // @[XRam.scala 144:57]
    end else begin
      reset_addr <= 10'h0; // @[XRam.scala 146:57]
    end
    REG <= io_addr_a; // @[XRam.scala 159:45]
    REG_1 <= io_addr_b; // @[XRam.scala 159:68]
    REG_2 <= io_wr_en_a; // @[XRam.scala 159:89]
    io_data_out_b_REG_max_field_num <= io_data_in_a_max_field_num; // @[XRam.scala 160:75]
    io_data_out_b_REG_field_type_0_is_repeated <= io_data_in_a_field_type_0_is_repeated; // @[XRam.scala 160:75]
    io_data_out_b_REG_field_type_0_field_type <= io_data_in_a_field_type_0_field_type; // @[XRam.scala 160:75]
    io_data_out_b_REG_field_type_0_sub_class_id <= io_data_in_a_field_type_0_sub_class_id; // @[XRam.scala 160:75]
    io_data_out_b_REG_field_type_1_is_repeated <= io_data_in_a_field_type_1_is_repeated; // @[XRam.scala 160:75]
    io_data_out_b_REG_field_type_1_field_type <= io_data_in_a_field_type_1_field_type; // @[XRam.scala 160:75]
    io_data_out_b_REG_field_type_1_sub_class_id <= io_data_in_a_field_type_1_sub_class_id; // @[XRam.scala 160:75]
    io_data_out_b_REG_field_type_2_is_repeated <= io_data_in_a_field_type_2_is_repeated; // @[XRam.scala 160:75]
    io_data_out_b_REG_field_type_2_field_type <= io_data_in_a_field_type_2_field_type; // @[XRam.scala 160:75]
    io_data_out_b_REG_field_type_2_sub_class_id <= io_data_in_a_field_type_2_sub_class_id; // @[XRam.scala 160:75]
    io_data_out_b_REG_field_type_3_is_repeated <= io_data_in_a_field_type_3_is_repeated; // @[XRam.scala 160:75]
    io_data_out_b_REG_field_type_3_field_type <= io_data_in_a_field_type_3_field_type; // @[XRam.scala 160:75]
    io_data_out_b_REG_field_type_3_sub_class_id <= io_data_in_a_field_type_3_sub_class_id; // @[XRam.scala 160:75]
    io_data_out_b_REG_field_type_4_is_repeated <= io_data_in_a_field_type_4_is_repeated; // @[XRam.scala 160:75]
    io_data_out_b_REG_field_type_4_field_type <= io_data_in_a_field_type_4_field_type; // @[XRam.scala 160:75]
    io_data_out_b_REG_field_type_4_sub_class_id <= io_data_in_a_field_type_4_sub_class_id; // @[XRam.scala 160:75]
    io_data_out_b_REG_field_type_5_is_repeated <= io_data_in_a_field_type_5_is_repeated; // @[XRam.scala 160:75]
    io_data_out_b_REG_field_type_5_field_type <= io_data_in_a_field_type_5_field_type; // @[XRam.scala 160:75]
    io_data_out_b_REG_field_type_5_sub_class_id <= io_data_in_a_field_type_5_sub_class_id; // @[XRam.scala 160:75]
    io_data_out_b_REG_field_type_6_is_repeated <= io_data_in_a_field_type_6_is_repeated; // @[XRam.scala 160:75]
    io_data_out_b_REG_field_type_6_field_type <= io_data_in_a_field_type_6_field_type; // @[XRam.scala 160:75]
    io_data_out_b_REG_field_type_6_sub_class_id <= io_data_in_a_field_type_6_sub_class_id; // @[XRam.scala 160:75]
    io_data_out_b_REG_field_type_7_is_repeated <= io_data_in_a_field_type_7_is_repeated; // @[XRam.scala 160:75]
    io_data_out_b_REG_field_type_7_field_type <= io_data_in_a_field_type_7_field_type; // @[XRam.scala 160:75]
    io_data_out_b_REG_field_type_7_sub_class_id <= io_data_in_a_field_type_7_sub_class_id; // @[XRam.scala 160:75]
    io_data_out_b_REG_field_type_8_is_repeated <= io_data_in_a_field_type_8_is_repeated; // @[XRam.scala 160:75]
    io_data_out_b_REG_field_type_8_field_type <= io_data_in_a_field_type_8_field_type; // @[XRam.scala 160:75]
    io_data_out_b_REG_field_type_8_sub_class_id <= io_data_in_a_field_type_8_sub_class_id; // @[XRam.scala 160:75]
    io_data_out_b_REG_field_type_9_is_repeated <= io_data_in_a_field_type_9_is_repeated; // @[XRam.scala 160:75]
    io_data_out_b_REG_field_type_9_field_type <= io_data_in_a_field_type_9_field_type; // @[XRam.scala 160:75]
    io_data_out_b_REG_field_type_9_sub_class_id <= io_data_in_a_field_type_9_sub_class_id; // @[XRam.scala 160:75]
    io_data_out_b_REG_field_type_10_is_repeated <= io_data_in_a_field_type_10_is_repeated; // @[XRam.scala 160:75]
    io_data_out_b_REG_field_type_10_field_type <= io_data_in_a_field_type_10_field_type; // @[XRam.scala 160:75]
    io_data_out_b_REG_field_type_10_sub_class_id <= io_data_in_a_field_type_10_sub_class_id; // @[XRam.scala 160:75]
    io_data_out_b_REG_field_type_11_is_repeated <= io_data_in_a_field_type_11_is_repeated; // @[XRam.scala 160:75]
    io_data_out_b_REG_field_type_11_field_type <= io_data_in_a_field_type_11_field_type; // @[XRam.scala 160:75]
    io_data_out_b_REG_field_type_11_sub_class_id <= io_data_in_a_field_type_11_sub_class_id; // @[XRam.scala 160:75]
    io_data_out_b_REG_field_type_12_is_repeated <= io_data_in_a_field_type_12_is_repeated; // @[XRam.scala 160:75]
    io_data_out_b_REG_field_type_12_field_type <= io_data_in_a_field_type_12_field_type; // @[XRam.scala 160:75]
    io_data_out_b_REG_field_type_12_sub_class_id <= io_data_in_a_field_type_12_sub_class_id; // @[XRam.scala 160:75]
    io_data_out_b_REG_field_type_13_is_repeated <= io_data_in_a_field_type_13_is_repeated; // @[XRam.scala 160:75]
    io_data_out_b_REG_field_type_13_field_type <= io_data_in_a_field_type_13_field_type; // @[XRam.scala 160:75]
    io_data_out_b_REG_field_type_13_sub_class_id <= io_data_in_a_field_type_13_sub_class_id; // @[XRam.scala 160:75]
    io_data_out_b_REG_field_type_14_is_repeated <= io_data_in_a_field_type_14_is_repeated; // @[XRam.scala 160:75]
    io_data_out_b_REG_field_type_14_field_type <= io_data_in_a_field_type_14_field_type; // @[XRam.scala 160:75]
    io_data_out_b_REG_field_type_14_sub_class_id <= io_data_in_a_field_type_14_sub_class_id; // @[XRam.scala 160:75]
    io_data_out_b_REG_field_type_15_is_repeated <= io_data_in_a_field_type_15_is_repeated; // @[XRam.scala 160:75]
    io_data_out_b_REG_field_type_15_field_type <= io_data_in_a_field_type_15_field_type; // @[XRam.scala 160:75]
    io_data_out_b_REG_field_type_15_sub_class_id <= io_data_in_a_field_type_15_sub_class_id; // @[XRam.scala 160:75]
    io_data_out_b_REG_field_type_16_is_repeated <= io_data_in_a_field_type_16_is_repeated; // @[XRam.scala 160:75]
    io_data_out_b_REG_field_type_16_field_type <= io_data_in_a_field_type_16_field_type; // @[XRam.scala 160:75]
    io_data_out_b_REG_field_type_16_sub_class_id <= io_data_in_a_field_type_16_sub_class_id; // @[XRam.scala 160:75]
    io_data_out_b_REG_field_type_17_is_repeated <= io_data_in_a_field_type_17_is_repeated; // @[XRam.scala 160:75]
    io_data_out_b_REG_field_type_17_field_type <= io_data_in_a_field_type_17_field_type; // @[XRam.scala 160:75]
    io_data_out_b_REG_field_type_17_sub_class_id <= io_data_in_a_field_type_17_sub_class_id; // @[XRam.scala 160:75]
    io_data_out_b_REG_field_type_18_is_repeated <= io_data_in_a_field_type_18_is_repeated; // @[XRam.scala 160:75]
    io_data_out_b_REG_field_type_18_field_type <= io_data_in_a_field_type_18_field_type; // @[XRam.scala 160:75]
    io_data_out_b_REG_field_type_18_sub_class_id <= io_data_in_a_field_type_18_sub_class_id; // @[XRam.scala 160:75]
    io_data_out_b_REG_field_type_19_is_repeated <= io_data_in_a_field_type_19_is_repeated; // @[XRam.scala 160:75]
    io_data_out_b_REG_field_type_19_field_type <= io_data_in_a_field_type_19_field_type; // @[XRam.scala 160:75]
    io_data_out_b_REG_field_type_19_sub_class_id <= io_data_in_a_field_type_19_sub_class_id; // @[XRam.scala 160:75]
    io_data_out_b_REG_field_type_20_is_repeated <= io_data_in_a_field_type_20_is_repeated; // @[XRam.scala 160:75]
    io_data_out_b_REG_field_type_20_field_type <= io_data_in_a_field_type_20_field_type; // @[XRam.scala 160:75]
    io_data_out_b_REG_field_type_20_sub_class_id <= io_data_in_a_field_type_20_sub_class_id; // @[XRam.scala 160:75]
    io_data_out_b_REG_field_type_21_is_repeated <= io_data_in_a_field_type_21_is_repeated; // @[XRam.scala 160:75]
    io_data_out_b_REG_field_type_21_field_type <= io_data_in_a_field_type_21_field_type; // @[XRam.scala 160:75]
    io_data_out_b_REG_field_type_21_sub_class_id <= io_data_in_a_field_type_21_sub_class_id; // @[XRam.scala 160:75]
    io_data_out_b_REG_field_type_22_is_repeated <= io_data_in_a_field_type_22_is_repeated; // @[XRam.scala 160:75]
    io_data_out_b_REG_field_type_22_field_type <= io_data_in_a_field_type_22_field_type; // @[XRam.scala 160:75]
    io_data_out_b_REG_field_type_22_sub_class_id <= io_data_in_a_field_type_22_sub_class_id; // @[XRam.scala 160:75]
    io_data_out_b_REG_field_type_23_is_repeated <= io_data_in_a_field_type_23_is_repeated; // @[XRam.scala 160:75]
    io_data_out_b_REG_field_type_23_field_type <= io_data_in_a_field_type_23_field_type; // @[XRam.scala 160:75]
    io_data_out_b_REG_field_type_23_sub_class_id <= io_data_in_a_field_type_23_sub_class_id; // @[XRam.scala 160:75]
    io_data_out_b_REG_field_type_24_is_repeated <= io_data_in_a_field_type_24_is_repeated; // @[XRam.scala 160:75]
    io_data_out_b_REG_field_type_24_field_type <= io_data_in_a_field_type_24_field_type; // @[XRam.scala 160:75]
    io_data_out_b_REG_field_type_24_sub_class_id <= io_data_in_a_field_type_24_sub_class_id; // @[XRam.scala 160:75]
    io_data_out_b_REG_field_type_25_is_repeated <= io_data_in_a_field_type_25_is_repeated; // @[XRam.scala 160:75]
    io_data_out_b_REG_field_type_25_field_type <= io_data_in_a_field_type_25_field_type; // @[XRam.scala 160:75]
    io_data_out_b_REG_field_type_25_sub_class_id <= io_data_in_a_field_type_25_sub_class_id; // @[XRam.scala 160:75]
    io_data_out_b_REG_field_type_26_is_repeated <= io_data_in_a_field_type_26_is_repeated; // @[XRam.scala 160:75]
    io_data_out_b_REG_field_type_26_field_type <= io_data_in_a_field_type_26_field_type; // @[XRam.scala 160:75]
    io_data_out_b_REG_field_type_26_sub_class_id <= io_data_in_a_field_type_26_sub_class_id; // @[XRam.scala 160:75]
    io_data_out_b_REG_field_type_27_is_repeated <= io_data_in_a_field_type_27_is_repeated; // @[XRam.scala 160:75]
    io_data_out_b_REG_field_type_27_field_type <= io_data_in_a_field_type_27_field_type; // @[XRam.scala 160:75]
    io_data_out_b_REG_field_type_27_sub_class_id <= io_data_in_a_field_type_27_sub_class_id; // @[XRam.scala 160:75]
    io_data_out_b_REG_field_type_28_is_repeated <= io_data_in_a_field_type_28_is_repeated; // @[XRam.scala 160:75]
    io_data_out_b_REG_field_type_28_field_type <= io_data_in_a_field_type_28_field_type; // @[XRam.scala 160:75]
    io_data_out_b_REG_field_type_28_sub_class_id <= io_data_in_a_field_type_28_sub_class_id; // @[XRam.scala 160:75]
    io_data_out_b_REG_field_type_29_is_repeated <= io_data_in_a_field_type_29_is_repeated; // @[XRam.scala 160:75]
    io_data_out_b_REG_field_type_29_field_type <= io_data_in_a_field_type_29_field_type; // @[XRam.scala 160:75]
    io_data_out_b_REG_field_type_29_sub_class_id <= io_data_in_a_field_type_29_sub_class_id; // @[XRam.scala 160:75]
    io_data_out_b_REG_field_type_30_is_repeated <= io_data_in_a_field_type_30_is_repeated; // @[XRam.scala 160:75]
    io_data_out_b_REG_field_type_30_field_type <= io_data_in_a_field_type_30_field_type; // @[XRam.scala 160:75]
    io_data_out_b_REG_field_type_30_sub_class_id <= io_data_in_a_field_type_30_sub_class_id; // @[XRam.scala 160:75]
    io_data_out_b_REG_field_type_31_is_repeated <= io_data_in_a_field_type_31_is_repeated; // @[XRam.scala 160:75]
    io_data_out_b_REG_field_type_31_field_type <= io_data_in_a_field_type_31_field_type; // @[XRam.scala 160:75]
    io_data_out_b_REG_field_type_31_sub_class_id <= io_data_in_a_field_type_31_sub_class_id; // @[XRam.scala 160:75]
    io_data_out_b_REG_field_type_32_is_repeated <= io_data_in_a_field_type_32_is_repeated; // @[XRam.scala 160:75]
    io_data_out_b_REG_field_type_32_field_type <= io_data_in_a_field_type_32_field_type; // @[XRam.scala 160:75]
    io_data_out_b_REG_field_type_32_sub_class_id <= io_data_in_a_field_type_32_sub_class_id; // @[XRam.scala 160:75]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  usr_rst_delay_r = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  usr_rst_delay_r_1 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  usr_rst_delay_r_2 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  usr_rst_delay = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  reset_addr = _RAND_4[9:0];
  _RAND_5 = {1{`RANDOM}};
  REG = _RAND_5[9:0];
  _RAND_6 = {1{`RANDOM}};
  REG_1 = _RAND_6[9:0];
  _RAND_7 = {1{`RANDOM}};
  REG_2 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  io_data_out_b_REG_max_field_num = _RAND_8[7:0];
  _RAND_9 = {1{`RANDOM}};
  io_data_out_b_REG_field_type_0_is_repeated = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  io_data_out_b_REG_field_type_0_field_type = _RAND_10[4:0];
  _RAND_11 = {1{`RANDOM}};
  io_data_out_b_REG_field_type_0_sub_class_id = _RAND_11[15:0];
  _RAND_12 = {1{`RANDOM}};
  io_data_out_b_REG_field_type_1_is_repeated = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  io_data_out_b_REG_field_type_1_field_type = _RAND_13[4:0];
  _RAND_14 = {1{`RANDOM}};
  io_data_out_b_REG_field_type_1_sub_class_id = _RAND_14[15:0];
  _RAND_15 = {1{`RANDOM}};
  io_data_out_b_REG_field_type_2_is_repeated = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  io_data_out_b_REG_field_type_2_field_type = _RAND_16[4:0];
  _RAND_17 = {1{`RANDOM}};
  io_data_out_b_REG_field_type_2_sub_class_id = _RAND_17[15:0];
  _RAND_18 = {1{`RANDOM}};
  io_data_out_b_REG_field_type_3_is_repeated = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  io_data_out_b_REG_field_type_3_field_type = _RAND_19[4:0];
  _RAND_20 = {1{`RANDOM}};
  io_data_out_b_REG_field_type_3_sub_class_id = _RAND_20[15:0];
  _RAND_21 = {1{`RANDOM}};
  io_data_out_b_REG_field_type_4_is_repeated = _RAND_21[0:0];
  _RAND_22 = {1{`RANDOM}};
  io_data_out_b_REG_field_type_4_field_type = _RAND_22[4:0];
  _RAND_23 = {1{`RANDOM}};
  io_data_out_b_REG_field_type_4_sub_class_id = _RAND_23[15:0];
  _RAND_24 = {1{`RANDOM}};
  io_data_out_b_REG_field_type_5_is_repeated = _RAND_24[0:0];
  _RAND_25 = {1{`RANDOM}};
  io_data_out_b_REG_field_type_5_field_type = _RAND_25[4:0];
  _RAND_26 = {1{`RANDOM}};
  io_data_out_b_REG_field_type_5_sub_class_id = _RAND_26[15:0];
  _RAND_27 = {1{`RANDOM}};
  io_data_out_b_REG_field_type_6_is_repeated = _RAND_27[0:0];
  _RAND_28 = {1{`RANDOM}};
  io_data_out_b_REG_field_type_6_field_type = _RAND_28[4:0];
  _RAND_29 = {1{`RANDOM}};
  io_data_out_b_REG_field_type_6_sub_class_id = _RAND_29[15:0];
  _RAND_30 = {1{`RANDOM}};
  io_data_out_b_REG_field_type_7_is_repeated = _RAND_30[0:0];
  _RAND_31 = {1{`RANDOM}};
  io_data_out_b_REG_field_type_7_field_type = _RAND_31[4:0];
  _RAND_32 = {1{`RANDOM}};
  io_data_out_b_REG_field_type_7_sub_class_id = _RAND_32[15:0];
  _RAND_33 = {1{`RANDOM}};
  io_data_out_b_REG_field_type_8_is_repeated = _RAND_33[0:0];
  _RAND_34 = {1{`RANDOM}};
  io_data_out_b_REG_field_type_8_field_type = _RAND_34[4:0];
  _RAND_35 = {1{`RANDOM}};
  io_data_out_b_REG_field_type_8_sub_class_id = _RAND_35[15:0];
  _RAND_36 = {1{`RANDOM}};
  io_data_out_b_REG_field_type_9_is_repeated = _RAND_36[0:0];
  _RAND_37 = {1{`RANDOM}};
  io_data_out_b_REG_field_type_9_field_type = _RAND_37[4:0];
  _RAND_38 = {1{`RANDOM}};
  io_data_out_b_REG_field_type_9_sub_class_id = _RAND_38[15:0];
  _RAND_39 = {1{`RANDOM}};
  io_data_out_b_REG_field_type_10_is_repeated = _RAND_39[0:0];
  _RAND_40 = {1{`RANDOM}};
  io_data_out_b_REG_field_type_10_field_type = _RAND_40[4:0];
  _RAND_41 = {1{`RANDOM}};
  io_data_out_b_REG_field_type_10_sub_class_id = _RAND_41[15:0];
  _RAND_42 = {1{`RANDOM}};
  io_data_out_b_REG_field_type_11_is_repeated = _RAND_42[0:0];
  _RAND_43 = {1{`RANDOM}};
  io_data_out_b_REG_field_type_11_field_type = _RAND_43[4:0];
  _RAND_44 = {1{`RANDOM}};
  io_data_out_b_REG_field_type_11_sub_class_id = _RAND_44[15:0];
  _RAND_45 = {1{`RANDOM}};
  io_data_out_b_REG_field_type_12_is_repeated = _RAND_45[0:0];
  _RAND_46 = {1{`RANDOM}};
  io_data_out_b_REG_field_type_12_field_type = _RAND_46[4:0];
  _RAND_47 = {1{`RANDOM}};
  io_data_out_b_REG_field_type_12_sub_class_id = _RAND_47[15:0];
  _RAND_48 = {1{`RANDOM}};
  io_data_out_b_REG_field_type_13_is_repeated = _RAND_48[0:0];
  _RAND_49 = {1{`RANDOM}};
  io_data_out_b_REG_field_type_13_field_type = _RAND_49[4:0];
  _RAND_50 = {1{`RANDOM}};
  io_data_out_b_REG_field_type_13_sub_class_id = _RAND_50[15:0];
  _RAND_51 = {1{`RANDOM}};
  io_data_out_b_REG_field_type_14_is_repeated = _RAND_51[0:0];
  _RAND_52 = {1{`RANDOM}};
  io_data_out_b_REG_field_type_14_field_type = _RAND_52[4:0];
  _RAND_53 = {1{`RANDOM}};
  io_data_out_b_REG_field_type_14_sub_class_id = _RAND_53[15:0];
  _RAND_54 = {1{`RANDOM}};
  io_data_out_b_REG_field_type_15_is_repeated = _RAND_54[0:0];
  _RAND_55 = {1{`RANDOM}};
  io_data_out_b_REG_field_type_15_field_type = _RAND_55[4:0];
  _RAND_56 = {1{`RANDOM}};
  io_data_out_b_REG_field_type_15_sub_class_id = _RAND_56[15:0];
  _RAND_57 = {1{`RANDOM}};
  io_data_out_b_REG_field_type_16_is_repeated = _RAND_57[0:0];
  _RAND_58 = {1{`RANDOM}};
  io_data_out_b_REG_field_type_16_field_type = _RAND_58[4:0];
  _RAND_59 = {1{`RANDOM}};
  io_data_out_b_REG_field_type_16_sub_class_id = _RAND_59[15:0];
  _RAND_60 = {1{`RANDOM}};
  io_data_out_b_REG_field_type_17_is_repeated = _RAND_60[0:0];
  _RAND_61 = {1{`RANDOM}};
  io_data_out_b_REG_field_type_17_field_type = _RAND_61[4:0];
  _RAND_62 = {1{`RANDOM}};
  io_data_out_b_REG_field_type_17_sub_class_id = _RAND_62[15:0];
  _RAND_63 = {1{`RANDOM}};
  io_data_out_b_REG_field_type_18_is_repeated = _RAND_63[0:0];
  _RAND_64 = {1{`RANDOM}};
  io_data_out_b_REG_field_type_18_field_type = _RAND_64[4:0];
  _RAND_65 = {1{`RANDOM}};
  io_data_out_b_REG_field_type_18_sub_class_id = _RAND_65[15:0];
  _RAND_66 = {1{`RANDOM}};
  io_data_out_b_REG_field_type_19_is_repeated = _RAND_66[0:0];
  _RAND_67 = {1{`RANDOM}};
  io_data_out_b_REG_field_type_19_field_type = _RAND_67[4:0];
  _RAND_68 = {1{`RANDOM}};
  io_data_out_b_REG_field_type_19_sub_class_id = _RAND_68[15:0];
  _RAND_69 = {1{`RANDOM}};
  io_data_out_b_REG_field_type_20_is_repeated = _RAND_69[0:0];
  _RAND_70 = {1{`RANDOM}};
  io_data_out_b_REG_field_type_20_field_type = _RAND_70[4:0];
  _RAND_71 = {1{`RANDOM}};
  io_data_out_b_REG_field_type_20_sub_class_id = _RAND_71[15:0];
  _RAND_72 = {1{`RANDOM}};
  io_data_out_b_REG_field_type_21_is_repeated = _RAND_72[0:0];
  _RAND_73 = {1{`RANDOM}};
  io_data_out_b_REG_field_type_21_field_type = _RAND_73[4:0];
  _RAND_74 = {1{`RANDOM}};
  io_data_out_b_REG_field_type_21_sub_class_id = _RAND_74[15:0];
  _RAND_75 = {1{`RANDOM}};
  io_data_out_b_REG_field_type_22_is_repeated = _RAND_75[0:0];
  _RAND_76 = {1{`RANDOM}};
  io_data_out_b_REG_field_type_22_field_type = _RAND_76[4:0];
  _RAND_77 = {1{`RANDOM}};
  io_data_out_b_REG_field_type_22_sub_class_id = _RAND_77[15:0];
  _RAND_78 = {1{`RANDOM}};
  io_data_out_b_REG_field_type_23_is_repeated = _RAND_78[0:0];
  _RAND_79 = {1{`RANDOM}};
  io_data_out_b_REG_field_type_23_field_type = _RAND_79[4:0];
  _RAND_80 = {1{`RANDOM}};
  io_data_out_b_REG_field_type_23_sub_class_id = _RAND_80[15:0];
  _RAND_81 = {1{`RANDOM}};
  io_data_out_b_REG_field_type_24_is_repeated = _RAND_81[0:0];
  _RAND_82 = {1{`RANDOM}};
  io_data_out_b_REG_field_type_24_field_type = _RAND_82[4:0];
  _RAND_83 = {1{`RANDOM}};
  io_data_out_b_REG_field_type_24_sub_class_id = _RAND_83[15:0];
  _RAND_84 = {1{`RANDOM}};
  io_data_out_b_REG_field_type_25_is_repeated = _RAND_84[0:0];
  _RAND_85 = {1{`RANDOM}};
  io_data_out_b_REG_field_type_25_field_type = _RAND_85[4:0];
  _RAND_86 = {1{`RANDOM}};
  io_data_out_b_REG_field_type_25_sub_class_id = _RAND_86[15:0];
  _RAND_87 = {1{`RANDOM}};
  io_data_out_b_REG_field_type_26_is_repeated = _RAND_87[0:0];
  _RAND_88 = {1{`RANDOM}};
  io_data_out_b_REG_field_type_26_field_type = _RAND_88[4:0];
  _RAND_89 = {1{`RANDOM}};
  io_data_out_b_REG_field_type_26_sub_class_id = _RAND_89[15:0];
  _RAND_90 = {1{`RANDOM}};
  io_data_out_b_REG_field_type_27_is_repeated = _RAND_90[0:0];
  _RAND_91 = {1{`RANDOM}};
  io_data_out_b_REG_field_type_27_field_type = _RAND_91[4:0];
  _RAND_92 = {1{`RANDOM}};
  io_data_out_b_REG_field_type_27_sub_class_id = _RAND_92[15:0];
  _RAND_93 = {1{`RANDOM}};
  io_data_out_b_REG_field_type_28_is_repeated = _RAND_93[0:0];
  _RAND_94 = {1{`RANDOM}};
  io_data_out_b_REG_field_type_28_field_type = _RAND_94[4:0];
  _RAND_95 = {1{`RANDOM}};
  io_data_out_b_REG_field_type_28_sub_class_id = _RAND_95[15:0];
  _RAND_96 = {1{`RANDOM}};
  io_data_out_b_REG_field_type_29_is_repeated = _RAND_96[0:0];
  _RAND_97 = {1{`RANDOM}};
  io_data_out_b_REG_field_type_29_field_type = _RAND_97[4:0];
  _RAND_98 = {1{`RANDOM}};
  io_data_out_b_REG_field_type_29_sub_class_id = _RAND_98[15:0];
  _RAND_99 = {1{`RANDOM}};
  io_data_out_b_REG_field_type_30_is_repeated = _RAND_99[0:0];
  _RAND_100 = {1{`RANDOM}};
  io_data_out_b_REG_field_type_30_field_type = _RAND_100[4:0];
  _RAND_101 = {1{`RANDOM}};
  io_data_out_b_REG_field_type_30_sub_class_id = _RAND_101[15:0];
  _RAND_102 = {1{`RANDOM}};
  io_data_out_b_REG_field_type_31_is_repeated = _RAND_102[0:0];
  _RAND_103 = {1{`RANDOM}};
  io_data_out_b_REG_field_type_31_field_type = _RAND_103[4:0];
  _RAND_104 = {1{`RANDOM}};
  io_data_out_b_REG_field_type_31_sub_class_id = _RAND_104[15:0];
  _RAND_105 = {1{`RANDOM}};
  io_data_out_b_REG_field_type_32_is_repeated = _RAND_105[0:0];
  _RAND_106 = {1{`RANDOM}};
  io_data_out_b_REG_field_type_32_field_type = _RAND_106[4:0];
  _RAND_107 = {1{`RANDOM}};
  io_data_out_b_REG_field_type_32_sub_class_id = _RAND_107[15:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ClassMetaTable(
  input         clock,
  input         reset,
  output        io_class_meta_init_ready,
  input         io_class_meta_init_valid,
  input  [9:0]  io_class_meta_init_bits_class_id,
  input  [15:0] io_class_meta_init_bits_desc_state_class_length,
  input  [7:0]  io_class_meta_init_bits_desc_state_max_field_num,
  input         io_class_meta_init_bits_desc_state_field_type_0_is_repeated,
  input  [4:0]  io_class_meta_init_bits_desc_state_field_type_0_field_type,
  input  [15:0] io_class_meta_init_bits_desc_state_field_type_0_sub_class_id,
  input         io_class_meta_init_bits_desc_state_field_type_0_is_host,
  input         io_class_meta_init_bits_desc_state_field_type_1_is_repeated,
  input  [4:0]  io_class_meta_init_bits_desc_state_field_type_1_field_type,
  input  [15:0] io_class_meta_init_bits_desc_state_field_type_1_sub_class_id,
  input         io_class_meta_init_bits_desc_state_field_type_1_is_host,
  input         io_class_meta_init_bits_desc_state_field_type_2_is_repeated,
  input  [4:0]  io_class_meta_init_bits_desc_state_field_type_2_field_type,
  input  [15:0] io_class_meta_init_bits_desc_state_field_type_2_sub_class_id,
  input         io_class_meta_init_bits_desc_state_field_type_2_is_host,
  input         io_class_meta_init_bits_desc_state_field_type_3_is_repeated,
  input  [4:0]  io_class_meta_init_bits_desc_state_field_type_3_field_type,
  input  [15:0] io_class_meta_init_bits_desc_state_field_type_3_sub_class_id,
  input         io_class_meta_init_bits_desc_state_field_type_3_is_host,
  input         io_class_meta_init_bits_desc_state_field_type_4_is_repeated,
  input  [4:0]  io_class_meta_init_bits_desc_state_field_type_4_field_type,
  input  [15:0] io_class_meta_init_bits_desc_state_field_type_4_sub_class_id,
  input         io_class_meta_init_bits_desc_state_field_type_4_is_host,
  input         io_class_meta_init_bits_desc_state_field_type_5_is_repeated,
  input  [4:0]  io_class_meta_init_bits_desc_state_field_type_5_field_type,
  input  [15:0] io_class_meta_init_bits_desc_state_field_type_5_sub_class_id,
  input         io_class_meta_init_bits_desc_state_field_type_5_is_host,
  input         io_class_meta_init_bits_desc_state_field_type_6_is_repeated,
  input  [4:0]  io_class_meta_init_bits_desc_state_field_type_6_field_type,
  input  [15:0] io_class_meta_init_bits_desc_state_field_type_6_sub_class_id,
  input         io_class_meta_init_bits_desc_state_field_type_6_is_host,
  input         io_class_meta_init_bits_desc_state_field_type_7_is_repeated,
  input  [4:0]  io_class_meta_init_bits_desc_state_field_type_7_field_type,
  input  [15:0] io_class_meta_init_bits_desc_state_field_type_7_sub_class_id,
  input         io_class_meta_init_bits_desc_state_field_type_7_is_host,
  input         io_class_meta_init_bits_desc_state_field_type_8_is_repeated,
  input  [4:0]  io_class_meta_init_bits_desc_state_field_type_8_field_type,
  input  [15:0] io_class_meta_init_bits_desc_state_field_type_8_sub_class_id,
  input         io_class_meta_init_bits_desc_state_field_type_8_is_host,
  input         io_class_meta_init_bits_desc_state_field_type_9_is_repeated,
  input  [4:0]  io_class_meta_init_bits_desc_state_field_type_9_field_type,
  input  [15:0] io_class_meta_init_bits_desc_state_field_type_9_sub_class_id,
  input         io_class_meta_init_bits_desc_state_field_type_9_is_host,
  input         io_class_meta_init_bits_desc_state_field_type_10_is_repeated,
  input  [4:0]  io_class_meta_init_bits_desc_state_field_type_10_field_type,
  input  [15:0] io_class_meta_init_bits_desc_state_field_type_10_sub_class_id,
  input         io_class_meta_init_bits_desc_state_field_type_10_is_host,
  input         io_class_meta_init_bits_desc_state_field_type_11_is_repeated,
  input  [4:0]  io_class_meta_init_bits_desc_state_field_type_11_field_type,
  input  [15:0] io_class_meta_init_bits_desc_state_field_type_11_sub_class_id,
  input         io_class_meta_init_bits_desc_state_field_type_11_is_host,
  input         io_class_meta_init_bits_desc_state_field_type_12_is_repeated,
  input  [4:0]  io_class_meta_init_bits_desc_state_field_type_12_field_type,
  input  [15:0] io_class_meta_init_bits_desc_state_field_type_12_sub_class_id,
  input         io_class_meta_init_bits_desc_state_field_type_12_is_host,
  input         io_class_meta_init_bits_desc_state_field_type_13_is_repeated,
  input  [4:0]  io_class_meta_init_bits_desc_state_field_type_13_field_type,
  input  [15:0] io_class_meta_init_bits_desc_state_field_type_13_sub_class_id,
  input         io_class_meta_init_bits_desc_state_field_type_13_is_host,
  input         io_class_meta_init_bits_desc_state_field_type_14_is_repeated,
  input  [4:0]  io_class_meta_init_bits_desc_state_field_type_14_field_type,
  input  [15:0] io_class_meta_init_bits_desc_state_field_type_14_sub_class_id,
  input         io_class_meta_init_bits_desc_state_field_type_14_is_host,
  input         io_class_meta_init_bits_desc_state_field_type_15_is_repeated,
  input  [4:0]  io_class_meta_init_bits_desc_state_field_type_15_field_type,
  input  [15:0] io_class_meta_init_bits_desc_state_field_type_15_sub_class_id,
  input         io_class_meta_init_bits_desc_state_field_type_15_is_host,
  input         io_class_meta_init_bits_desc_state_field_type_16_is_repeated,
  input  [4:0]  io_class_meta_init_bits_desc_state_field_type_16_field_type,
  input  [15:0] io_class_meta_init_bits_desc_state_field_type_16_sub_class_id,
  input         io_class_meta_init_bits_desc_state_field_type_16_is_host,
  input         io_class_meta_init_bits_desc_state_field_type_17_is_repeated,
  input  [4:0]  io_class_meta_init_bits_desc_state_field_type_17_field_type,
  input  [15:0] io_class_meta_init_bits_desc_state_field_type_17_sub_class_id,
  input         io_class_meta_init_bits_desc_state_field_type_17_is_host,
  input         io_class_meta_init_bits_desc_state_field_type_18_is_repeated,
  input  [4:0]  io_class_meta_init_bits_desc_state_field_type_18_field_type,
  input  [15:0] io_class_meta_init_bits_desc_state_field_type_18_sub_class_id,
  input         io_class_meta_init_bits_desc_state_field_type_18_is_host,
  input         io_class_meta_init_bits_desc_state_field_type_19_is_repeated,
  input  [4:0]  io_class_meta_init_bits_desc_state_field_type_19_field_type,
  input  [15:0] io_class_meta_init_bits_desc_state_field_type_19_sub_class_id,
  input         io_class_meta_init_bits_desc_state_field_type_19_is_host,
  input         io_class_meta_init_bits_desc_state_field_type_20_is_repeated,
  input  [4:0]  io_class_meta_init_bits_desc_state_field_type_20_field_type,
  input  [15:0] io_class_meta_init_bits_desc_state_field_type_20_sub_class_id,
  input         io_class_meta_init_bits_desc_state_field_type_20_is_host,
  input         io_class_meta_init_bits_desc_state_field_type_21_is_repeated,
  input  [4:0]  io_class_meta_init_bits_desc_state_field_type_21_field_type,
  input  [15:0] io_class_meta_init_bits_desc_state_field_type_21_sub_class_id,
  input         io_class_meta_init_bits_desc_state_field_type_21_is_host,
  input         io_class_meta_init_bits_desc_state_field_type_22_is_repeated,
  input  [4:0]  io_class_meta_init_bits_desc_state_field_type_22_field_type,
  input  [15:0] io_class_meta_init_bits_desc_state_field_type_22_sub_class_id,
  input         io_class_meta_init_bits_desc_state_field_type_22_is_host,
  input         io_class_meta_init_bits_desc_state_field_type_23_is_repeated,
  input  [4:0]  io_class_meta_init_bits_desc_state_field_type_23_field_type,
  input  [15:0] io_class_meta_init_bits_desc_state_field_type_23_sub_class_id,
  input         io_class_meta_init_bits_desc_state_field_type_23_is_host,
  input         io_class_meta_init_bits_desc_state_field_type_24_is_repeated,
  input  [4:0]  io_class_meta_init_bits_desc_state_field_type_24_field_type,
  input  [15:0] io_class_meta_init_bits_desc_state_field_type_24_sub_class_id,
  input         io_class_meta_init_bits_desc_state_field_type_24_is_host,
  input         io_class_meta_init_bits_desc_state_field_type_25_is_repeated,
  input  [4:0]  io_class_meta_init_bits_desc_state_field_type_25_field_type,
  input  [15:0] io_class_meta_init_bits_desc_state_field_type_25_sub_class_id,
  input         io_class_meta_init_bits_desc_state_field_type_25_is_host,
  input         io_class_meta_init_bits_desc_state_field_type_26_is_repeated,
  input  [4:0]  io_class_meta_init_bits_desc_state_field_type_26_field_type,
  input  [15:0] io_class_meta_init_bits_desc_state_field_type_26_sub_class_id,
  input         io_class_meta_init_bits_desc_state_field_type_26_is_host,
  input         io_class_meta_init_bits_desc_state_field_type_27_is_repeated,
  input  [4:0]  io_class_meta_init_bits_desc_state_field_type_27_field_type,
  input  [15:0] io_class_meta_init_bits_desc_state_field_type_27_sub_class_id,
  input         io_class_meta_init_bits_desc_state_field_type_27_is_host,
  input         io_class_meta_init_bits_desc_state_field_type_28_is_repeated,
  input  [4:0]  io_class_meta_init_bits_desc_state_field_type_28_field_type,
  input  [15:0] io_class_meta_init_bits_desc_state_field_type_28_sub_class_id,
  input         io_class_meta_init_bits_desc_state_field_type_28_is_host,
  input         io_class_meta_init_bits_desc_state_field_type_29_is_repeated,
  input  [4:0]  io_class_meta_init_bits_desc_state_field_type_29_field_type,
  input  [15:0] io_class_meta_init_bits_desc_state_field_type_29_sub_class_id,
  input         io_class_meta_init_bits_desc_state_field_type_29_is_host,
  input         io_class_meta_init_bits_desc_state_field_type_30_is_repeated,
  input  [4:0]  io_class_meta_init_bits_desc_state_field_type_30_field_type,
  input  [15:0] io_class_meta_init_bits_desc_state_field_type_30_sub_class_id,
  input         io_class_meta_init_bits_desc_state_field_type_30_is_host,
  input         io_class_meta_init_bits_desc_state_field_type_31_is_repeated,
  input  [4:0]  io_class_meta_init_bits_desc_state_field_type_31_field_type,
  input  [15:0] io_class_meta_init_bits_desc_state_field_type_31_sub_class_id,
  input         io_class_meta_init_bits_desc_state_field_type_31_is_host,
  input         io_class_meta_init_bits_desc_state_field_type_32_is_repeated,
  input  [4:0]  io_class_meta_init_bits_desc_state_field_type_32_field_type,
  input  [15:0] io_class_meta_init_bits_desc_state_field_type_32_sub_class_id,
  input         io_class_meta_init_bits_desc_state_field_type_32_is_host,
  output        io_s_class_meta_req_ready,
  input         io_s_class_meta_req_valid,
  input  [9:0]  io_s_class_meta_req_bits_class_id,
  output        io_s_class_meta_rsp_valid,
  output [7:0]  io_s_class_meta_rsp_bits_class_meta_max_field_num,
  output        io_s_class_meta_rsp_bits_class_meta_field_type_0_is_repeated,
  output [4:0]  io_s_class_meta_rsp_bits_class_meta_field_type_0_field_type,
  output [15:0] io_s_class_meta_rsp_bits_class_meta_field_type_0_sub_class_id,
  output        io_s_class_meta_rsp_bits_class_meta_field_type_1_is_repeated,
  output [4:0]  io_s_class_meta_rsp_bits_class_meta_field_type_1_field_type,
  output [15:0] io_s_class_meta_rsp_bits_class_meta_field_type_1_sub_class_id,
  output        io_s_class_meta_rsp_bits_class_meta_field_type_2_is_repeated,
  output [4:0]  io_s_class_meta_rsp_bits_class_meta_field_type_2_field_type,
  output [15:0] io_s_class_meta_rsp_bits_class_meta_field_type_2_sub_class_id,
  output        io_s_class_meta_rsp_bits_class_meta_field_type_3_is_repeated,
  output [4:0]  io_s_class_meta_rsp_bits_class_meta_field_type_3_field_type,
  output [15:0] io_s_class_meta_rsp_bits_class_meta_field_type_3_sub_class_id,
  output        io_s_class_meta_rsp_bits_class_meta_field_type_4_is_repeated,
  output [4:0]  io_s_class_meta_rsp_bits_class_meta_field_type_4_field_type,
  output [15:0] io_s_class_meta_rsp_bits_class_meta_field_type_4_sub_class_id,
  output        io_s_class_meta_rsp_bits_class_meta_field_type_5_is_repeated,
  output [4:0]  io_s_class_meta_rsp_bits_class_meta_field_type_5_field_type,
  output [15:0] io_s_class_meta_rsp_bits_class_meta_field_type_5_sub_class_id,
  output        io_s_class_meta_rsp_bits_class_meta_field_type_6_is_repeated,
  output [4:0]  io_s_class_meta_rsp_bits_class_meta_field_type_6_field_type,
  output [15:0] io_s_class_meta_rsp_bits_class_meta_field_type_6_sub_class_id,
  output        io_s_class_meta_rsp_bits_class_meta_field_type_7_is_repeated,
  output [4:0]  io_s_class_meta_rsp_bits_class_meta_field_type_7_field_type,
  output [15:0] io_s_class_meta_rsp_bits_class_meta_field_type_7_sub_class_id,
  output        io_s_class_meta_rsp_bits_class_meta_field_type_8_is_repeated,
  output [4:0]  io_s_class_meta_rsp_bits_class_meta_field_type_8_field_type,
  output [15:0] io_s_class_meta_rsp_bits_class_meta_field_type_8_sub_class_id,
  output        io_s_class_meta_rsp_bits_class_meta_field_type_9_is_repeated,
  output [4:0]  io_s_class_meta_rsp_bits_class_meta_field_type_9_field_type,
  output [15:0] io_s_class_meta_rsp_bits_class_meta_field_type_9_sub_class_id,
  output        io_s_class_meta_rsp_bits_class_meta_field_type_10_is_repeated,
  output [4:0]  io_s_class_meta_rsp_bits_class_meta_field_type_10_field_type,
  output [15:0] io_s_class_meta_rsp_bits_class_meta_field_type_10_sub_class_id,
  output        io_s_class_meta_rsp_bits_class_meta_field_type_11_is_repeated,
  output [4:0]  io_s_class_meta_rsp_bits_class_meta_field_type_11_field_type,
  output [15:0] io_s_class_meta_rsp_bits_class_meta_field_type_11_sub_class_id,
  output        io_s_class_meta_rsp_bits_class_meta_field_type_12_is_repeated,
  output [4:0]  io_s_class_meta_rsp_bits_class_meta_field_type_12_field_type,
  output [15:0] io_s_class_meta_rsp_bits_class_meta_field_type_12_sub_class_id,
  output        io_s_class_meta_rsp_bits_class_meta_field_type_13_is_repeated,
  output [4:0]  io_s_class_meta_rsp_bits_class_meta_field_type_13_field_type,
  output [15:0] io_s_class_meta_rsp_bits_class_meta_field_type_13_sub_class_id,
  output        io_s_class_meta_rsp_bits_class_meta_field_type_14_is_repeated,
  output [4:0]  io_s_class_meta_rsp_bits_class_meta_field_type_14_field_type,
  output [15:0] io_s_class_meta_rsp_bits_class_meta_field_type_14_sub_class_id,
  output        io_s_class_meta_rsp_bits_class_meta_field_type_15_is_repeated,
  output [4:0]  io_s_class_meta_rsp_bits_class_meta_field_type_15_field_type,
  output [15:0] io_s_class_meta_rsp_bits_class_meta_field_type_15_sub_class_id,
  output        io_s_class_meta_rsp_bits_class_meta_field_type_16_is_repeated,
  output [4:0]  io_s_class_meta_rsp_bits_class_meta_field_type_16_field_type,
  output [15:0] io_s_class_meta_rsp_bits_class_meta_field_type_16_sub_class_id,
  output        io_s_class_meta_rsp_bits_class_meta_field_type_17_is_repeated,
  output [4:0]  io_s_class_meta_rsp_bits_class_meta_field_type_17_field_type,
  output [15:0] io_s_class_meta_rsp_bits_class_meta_field_type_17_sub_class_id,
  output        io_s_class_meta_rsp_bits_class_meta_field_type_18_is_repeated,
  output [4:0]  io_s_class_meta_rsp_bits_class_meta_field_type_18_field_type,
  output [15:0] io_s_class_meta_rsp_bits_class_meta_field_type_18_sub_class_id,
  output        io_s_class_meta_rsp_bits_class_meta_field_type_19_is_repeated,
  output [4:0]  io_s_class_meta_rsp_bits_class_meta_field_type_19_field_type,
  output [15:0] io_s_class_meta_rsp_bits_class_meta_field_type_19_sub_class_id,
  output        io_s_class_meta_rsp_bits_class_meta_field_type_20_is_repeated,
  output [4:0]  io_s_class_meta_rsp_bits_class_meta_field_type_20_field_type,
  output [15:0] io_s_class_meta_rsp_bits_class_meta_field_type_20_sub_class_id,
  output        io_s_class_meta_rsp_bits_class_meta_field_type_21_is_repeated,
  output [4:0]  io_s_class_meta_rsp_bits_class_meta_field_type_21_field_type,
  output [15:0] io_s_class_meta_rsp_bits_class_meta_field_type_21_sub_class_id,
  output        io_s_class_meta_rsp_bits_class_meta_field_type_22_is_repeated,
  output [4:0]  io_s_class_meta_rsp_bits_class_meta_field_type_22_field_type,
  output [15:0] io_s_class_meta_rsp_bits_class_meta_field_type_22_sub_class_id,
  output        io_s_class_meta_rsp_bits_class_meta_field_type_23_is_repeated,
  output [4:0]  io_s_class_meta_rsp_bits_class_meta_field_type_23_field_type,
  output [15:0] io_s_class_meta_rsp_bits_class_meta_field_type_23_sub_class_id,
  output        io_s_class_meta_rsp_bits_class_meta_field_type_24_is_repeated,
  output [4:0]  io_s_class_meta_rsp_bits_class_meta_field_type_24_field_type,
  output [15:0] io_s_class_meta_rsp_bits_class_meta_field_type_24_sub_class_id,
  output        io_s_class_meta_rsp_bits_class_meta_field_type_25_is_repeated,
  output [4:0]  io_s_class_meta_rsp_bits_class_meta_field_type_25_field_type,
  output [15:0] io_s_class_meta_rsp_bits_class_meta_field_type_25_sub_class_id,
  output        io_s_class_meta_rsp_bits_class_meta_field_type_26_is_repeated,
  output [4:0]  io_s_class_meta_rsp_bits_class_meta_field_type_26_field_type,
  output [15:0] io_s_class_meta_rsp_bits_class_meta_field_type_26_sub_class_id,
  output        io_s_class_meta_rsp_bits_class_meta_field_type_27_is_repeated,
  output [4:0]  io_s_class_meta_rsp_bits_class_meta_field_type_27_field_type,
  output [15:0] io_s_class_meta_rsp_bits_class_meta_field_type_27_sub_class_id,
  output        io_s_class_meta_rsp_bits_class_meta_field_type_28_is_repeated,
  output [4:0]  io_s_class_meta_rsp_bits_class_meta_field_type_28_field_type,
  output [15:0] io_s_class_meta_rsp_bits_class_meta_field_type_28_sub_class_id,
  output        io_s_class_meta_rsp_bits_class_meta_field_type_29_is_repeated,
  output [4:0]  io_s_class_meta_rsp_bits_class_meta_field_type_29_field_type,
  output [15:0] io_s_class_meta_rsp_bits_class_meta_field_type_29_sub_class_id,
  output        io_s_class_meta_rsp_bits_class_meta_field_type_30_is_repeated,
  output [4:0]  io_s_class_meta_rsp_bits_class_meta_field_type_30_field_type,
  output [15:0] io_s_class_meta_rsp_bits_class_meta_field_type_30_sub_class_id,
  output        io_s_class_meta_rsp_bits_class_meta_field_type_31_is_repeated,
  output [4:0]  io_s_class_meta_rsp_bits_class_meta_field_type_31_field_type,
  output [15:0] io_s_class_meta_rsp_bits_class_meta_field_type_31_sub_class_id,
  output        io_s_class_meta_rsp_bits_class_meta_field_type_32_is_repeated,
  output [4:0]  io_s_class_meta_rsp_bits_class_meta_field_type_32_field_type,
  output [15:0] io_s_class_meta_rsp_bits_class_meta_field_type_32_sub_class_id,
  output [31:0] counter_5
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  wire  s_class_meta_req_fifo_clock; // @[XQueue.scala 35:23]
  wire  s_class_meta_req_fifo_reset; // @[XQueue.scala 35:23]
  wire  s_class_meta_req_fifo_io_in_ready; // @[XQueue.scala 35:23]
  wire  s_class_meta_req_fifo_io_in_valid; // @[XQueue.scala 35:23]
  wire [9:0] s_class_meta_req_fifo_io_in_bits_class_id; // @[XQueue.scala 35:23]
  wire  s_class_meta_req_fifo_io_out_ready; // @[XQueue.scala 35:23]
  wire  s_class_meta_req_fifo_io_out_valid; // @[XQueue.scala 35:23]
  wire [9:0] s_class_meta_req_fifo_io_out_bits_class_id; // @[XQueue.scala 35:23]
  wire  d_class_meta_req_fifo_clock; // @[XQueue.scala 35:23]
  wire  d_class_meta_req_fifo_reset; // @[XQueue.scala 35:23]
  wire  d_class_meta_req_fifo_io_in_ready; // @[XQueue.scala 35:23]
  wire  d_class_meta_req_fifo_io_in_valid; // @[XQueue.scala 35:23]
  wire [9:0] d_class_meta_req_fifo_io_in_bits_class_id; // @[XQueue.scala 35:23]
  wire  d_class_meta_req_fifo_io_out_ready; // @[XQueue.scala 35:23]
  wire  d_class_meta_req_fifo_io_out_valid; // @[XQueue.scala 35:23]
  wire [9:0] d_class_meta_req_fifo_io_out_bits_class_id; // @[XQueue.scala 35:23]
  wire  meta_table_clock; // @[XRam.scala 102:23]
  wire  meta_table_reset; // @[XRam.scala 102:23]
  wire [9:0] meta_table_io_addr_a; // @[XRam.scala 102:23]
  wire [9:0] meta_table_io_addr_b; // @[XRam.scala 102:23]
  wire  meta_table_io_wr_en_a; // @[XRam.scala 102:23]
  wire [15:0] meta_table_io_data_in_a_class_length; // @[XRam.scala 102:23]
  wire [7:0] meta_table_io_data_in_a_max_field_num; // @[XRam.scala 102:23]
  wire  meta_table_io_data_in_a_field_type_0_is_repeated; // @[XRam.scala 102:23]
  wire [4:0] meta_table_io_data_in_a_field_type_0_field_type; // @[XRam.scala 102:23]
  wire [15:0] meta_table_io_data_in_a_field_type_0_sub_class_id; // @[XRam.scala 102:23]
  wire  meta_table_io_data_in_a_field_type_0_is_host; // @[XRam.scala 102:23]
  wire  meta_table_io_data_in_a_field_type_1_is_repeated; // @[XRam.scala 102:23]
  wire [4:0] meta_table_io_data_in_a_field_type_1_field_type; // @[XRam.scala 102:23]
  wire [15:0] meta_table_io_data_in_a_field_type_1_sub_class_id; // @[XRam.scala 102:23]
  wire  meta_table_io_data_in_a_field_type_1_is_host; // @[XRam.scala 102:23]
  wire  meta_table_io_data_in_a_field_type_2_is_repeated; // @[XRam.scala 102:23]
  wire [4:0] meta_table_io_data_in_a_field_type_2_field_type; // @[XRam.scala 102:23]
  wire [15:0] meta_table_io_data_in_a_field_type_2_sub_class_id; // @[XRam.scala 102:23]
  wire  meta_table_io_data_in_a_field_type_2_is_host; // @[XRam.scala 102:23]
  wire  meta_table_io_data_in_a_field_type_3_is_repeated; // @[XRam.scala 102:23]
  wire [4:0] meta_table_io_data_in_a_field_type_3_field_type; // @[XRam.scala 102:23]
  wire [15:0] meta_table_io_data_in_a_field_type_3_sub_class_id; // @[XRam.scala 102:23]
  wire  meta_table_io_data_in_a_field_type_3_is_host; // @[XRam.scala 102:23]
  wire  meta_table_io_data_in_a_field_type_4_is_repeated; // @[XRam.scala 102:23]
  wire [4:0] meta_table_io_data_in_a_field_type_4_field_type; // @[XRam.scala 102:23]
  wire [15:0] meta_table_io_data_in_a_field_type_4_sub_class_id; // @[XRam.scala 102:23]
  wire  meta_table_io_data_in_a_field_type_4_is_host; // @[XRam.scala 102:23]
  wire  meta_table_io_data_in_a_field_type_5_is_repeated; // @[XRam.scala 102:23]
  wire [4:0] meta_table_io_data_in_a_field_type_5_field_type; // @[XRam.scala 102:23]
  wire [15:0] meta_table_io_data_in_a_field_type_5_sub_class_id; // @[XRam.scala 102:23]
  wire  meta_table_io_data_in_a_field_type_5_is_host; // @[XRam.scala 102:23]
  wire  meta_table_io_data_in_a_field_type_6_is_repeated; // @[XRam.scala 102:23]
  wire [4:0] meta_table_io_data_in_a_field_type_6_field_type; // @[XRam.scala 102:23]
  wire [15:0] meta_table_io_data_in_a_field_type_6_sub_class_id; // @[XRam.scala 102:23]
  wire  meta_table_io_data_in_a_field_type_6_is_host; // @[XRam.scala 102:23]
  wire  meta_table_io_data_in_a_field_type_7_is_repeated; // @[XRam.scala 102:23]
  wire [4:0] meta_table_io_data_in_a_field_type_7_field_type; // @[XRam.scala 102:23]
  wire [15:0] meta_table_io_data_in_a_field_type_7_sub_class_id; // @[XRam.scala 102:23]
  wire  meta_table_io_data_in_a_field_type_7_is_host; // @[XRam.scala 102:23]
  wire  meta_table_io_data_in_a_field_type_8_is_repeated; // @[XRam.scala 102:23]
  wire [4:0] meta_table_io_data_in_a_field_type_8_field_type; // @[XRam.scala 102:23]
  wire [15:0] meta_table_io_data_in_a_field_type_8_sub_class_id; // @[XRam.scala 102:23]
  wire  meta_table_io_data_in_a_field_type_8_is_host; // @[XRam.scala 102:23]
  wire  meta_table_io_data_in_a_field_type_9_is_repeated; // @[XRam.scala 102:23]
  wire [4:0] meta_table_io_data_in_a_field_type_9_field_type; // @[XRam.scala 102:23]
  wire [15:0] meta_table_io_data_in_a_field_type_9_sub_class_id; // @[XRam.scala 102:23]
  wire  meta_table_io_data_in_a_field_type_9_is_host; // @[XRam.scala 102:23]
  wire  meta_table_io_data_in_a_field_type_10_is_repeated; // @[XRam.scala 102:23]
  wire [4:0] meta_table_io_data_in_a_field_type_10_field_type; // @[XRam.scala 102:23]
  wire [15:0] meta_table_io_data_in_a_field_type_10_sub_class_id; // @[XRam.scala 102:23]
  wire  meta_table_io_data_in_a_field_type_10_is_host; // @[XRam.scala 102:23]
  wire  meta_table_io_data_in_a_field_type_11_is_repeated; // @[XRam.scala 102:23]
  wire [4:0] meta_table_io_data_in_a_field_type_11_field_type; // @[XRam.scala 102:23]
  wire [15:0] meta_table_io_data_in_a_field_type_11_sub_class_id; // @[XRam.scala 102:23]
  wire  meta_table_io_data_in_a_field_type_11_is_host; // @[XRam.scala 102:23]
  wire  meta_table_io_data_in_a_field_type_12_is_repeated; // @[XRam.scala 102:23]
  wire [4:0] meta_table_io_data_in_a_field_type_12_field_type; // @[XRam.scala 102:23]
  wire [15:0] meta_table_io_data_in_a_field_type_12_sub_class_id; // @[XRam.scala 102:23]
  wire  meta_table_io_data_in_a_field_type_12_is_host; // @[XRam.scala 102:23]
  wire  meta_table_io_data_in_a_field_type_13_is_repeated; // @[XRam.scala 102:23]
  wire [4:0] meta_table_io_data_in_a_field_type_13_field_type; // @[XRam.scala 102:23]
  wire [15:0] meta_table_io_data_in_a_field_type_13_sub_class_id; // @[XRam.scala 102:23]
  wire  meta_table_io_data_in_a_field_type_13_is_host; // @[XRam.scala 102:23]
  wire  meta_table_io_data_in_a_field_type_14_is_repeated; // @[XRam.scala 102:23]
  wire [4:0] meta_table_io_data_in_a_field_type_14_field_type; // @[XRam.scala 102:23]
  wire [15:0] meta_table_io_data_in_a_field_type_14_sub_class_id; // @[XRam.scala 102:23]
  wire  meta_table_io_data_in_a_field_type_14_is_host; // @[XRam.scala 102:23]
  wire  meta_table_io_data_in_a_field_type_15_is_repeated; // @[XRam.scala 102:23]
  wire [4:0] meta_table_io_data_in_a_field_type_15_field_type; // @[XRam.scala 102:23]
  wire [15:0] meta_table_io_data_in_a_field_type_15_sub_class_id; // @[XRam.scala 102:23]
  wire  meta_table_io_data_in_a_field_type_15_is_host; // @[XRam.scala 102:23]
  wire  meta_table_io_data_in_a_field_type_16_is_repeated; // @[XRam.scala 102:23]
  wire [4:0] meta_table_io_data_in_a_field_type_16_field_type; // @[XRam.scala 102:23]
  wire [15:0] meta_table_io_data_in_a_field_type_16_sub_class_id; // @[XRam.scala 102:23]
  wire  meta_table_io_data_in_a_field_type_16_is_host; // @[XRam.scala 102:23]
  wire  meta_table_io_data_in_a_field_type_17_is_repeated; // @[XRam.scala 102:23]
  wire [4:0] meta_table_io_data_in_a_field_type_17_field_type; // @[XRam.scala 102:23]
  wire [15:0] meta_table_io_data_in_a_field_type_17_sub_class_id; // @[XRam.scala 102:23]
  wire  meta_table_io_data_in_a_field_type_17_is_host; // @[XRam.scala 102:23]
  wire  meta_table_io_data_in_a_field_type_18_is_repeated; // @[XRam.scala 102:23]
  wire [4:0] meta_table_io_data_in_a_field_type_18_field_type; // @[XRam.scala 102:23]
  wire [15:0] meta_table_io_data_in_a_field_type_18_sub_class_id; // @[XRam.scala 102:23]
  wire  meta_table_io_data_in_a_field_type_18_is_host; // @[XRam.scala 102:23]
  wire  meta_table_io_data_in_a_field_type_19_is_repeated; // @[XRam.scala 102:23]
  wire [4:0] meta_table_io_data_in_a_field_type_19_field_type; // @[XRam.scala 102:23]
  wire [15:0] meta_table_io_data_in_a_field_type_19_sub_class_id; // @[XRam.scala 102:23]
  wire  meta_table_io_data_in_a_field_type_19_is_host; // @[XRam.scala 102:23]
  wire  meta_table_io_data_in_a_field_type_20_is_repeated; // @[XRam.scala 102:23]
  wire [4:0] meta_table_io_data_in_a_field_type_20_field_type; // @[XRam.scala 102:23]
  wire [15:0] meta_table_io_data_in_a_field_type_20_sub_class_id; // @[XRam.scala 102:23]
  wire  meta_table_io_data_in_a_field_type_20_is_host; // @[XRam.scala 102:23]
  wire  meta_table_io_data_in_a_field_type_21_is_repeated; // @[XRam.scala 102:23]
  wire [4:0] meta_table_io_data_in_a_field_type_21_field_type; // @[XRam.scala 102:23]
  wire [15:0] meta_table_io_data_in_a_field_type_21_sub_class_id; // @[XRam.scala 102:23]
  wire  meta_table_io_data_in_a_field_type_21_is_host; // @[XRam.scala 102:23]
  wire  meta_table_io_data_in_a_field_type_22_is_repeated; // @[XRam.scala 102:23]
  wire [4:0] meta_table_io_data_in_a_field_type_22_field_type; // @[XRam.scala 102:23]
  wire [15:0] meta_table_io_data_in_a_field_type_22_sub_class_id; // @[XRam.scala 102:23]
  wire  meta_table_io_data_in_a_field_type_22_is_host; // @[XRam.scala 102:23]
  wire  meta_table_io_data_in_a_field_type_23_is_repeated; // @[XRam.scala 102:23]
  wire [4:0] meta_table_io_data_in_a_field_type_23_field_type; // @[XRam.scala 102:23]
  wire [15:0] meta_table_io_data_in_a_field_type_23_sub_class_id; // @[XRam.scala 102:23]
  wire  meta_table_io_data_in_a_field_type_23_is_host; // @[XRam.scala 102:23]
  wire  meta_table_io_data_in_a_field_type_24_is_repeated; // @[XRam.scala 102:23]
  wire [4:0] meta_table_io_data_in_a_field_type_24_field_type; // @[XRam.scala 102:23]
  wire [15:0] meta_table_io_data_in_a_field_type_24_sub_class_id; // @[XRam.scala 102:23]
  wire  meta_table_io_data_in_a_field_type_24_is_host; // @[XRam.scala 102:23]
  wire  meta_table_io_data_in_a_field_type_25_is_repeated; // @[XRam.scala 102:23]
  wire [4:0] meta_table_io_data_in_a_field_type_25_field_type; // @[XRam.scala 102:23]
  wire [15:0] meta_table_io_data_in_a_field_type_25_sub_class_id; // @[XRam.scala 102:23]
  wire  meta_table_io_data_in_a_field_type_25_is_host; // @[XRam.scala 102:23]
  wire  meta_table_io_data_in_a_field_type_26_is_repeated; // @[XRam.scala 102:23]
  wire [4:0] meta_table_io_data_in_a_field_type_26_field_type; // @[XRam.scala 102:23]
  wire [15:0] meta_table_io_data_in_a_field_type_26_sub_class_id; // @[XRam.scala 102:23]
  wire  meta_table_io_data_in_a_field_type_26_is_host; // @[XRam.scala 102:23]
  wire  meta_table_io_data_in_a_field_type_27_is_repeated; // @[XRam.scala 102:23]
  wire [4:0] meta_table_io_data_in_a_field_type_27_field_type; // @[XRam.scala 102:23]
  wire [15:0] meta_table_io_data_in_a_field_type_27_sub_class_id; // @[XRam.scala 102:23]
  wire  meta_table_io_data_in_a_field_type_27_is_host; // @[XRam.scala 102:23]
  wire  meta_table_io_data_in_a_field_type_28_is_repeated; // @[XRam.scala 102:23]
  wire [4:0] meta_table_io_data_in_a_field_type_28_field_type; // @[XRam.scala 102:23]
  wire [15:0] meta_table_io_data_in_a_field_type_28_sub_class_id; // @[XRam.scala 102:23]
  wire  meta_table_io_data_in_a_field_type_28_is_host; // @[XRam.scala 102:23]
  wire  meta_table_io_data_in_a_field_type_29_is_repeated; // @[XRam.scala 102:23]
  wire [4:0] meta_table_io_data_in_a_field_type_29_field_type; // @[XRam.scala 102:23]
  wire [15:0] meta_table_io_data_in_a_field_type_29_sub_class_id; // @[XRam.scala 102:23]
  wire  meta_table_io_data_in_a_field_type_29_is_host; // @[XRam.scala 102:23]
  wire  meta_table_io_data_in_a_field_type_30_is_repeated; // @[XRam.scala 102:23]
  wire [4:0] meta_table_io_data_in_a_field_type_30_field_type; // @[XRam.scala 102:23]
  wire [15:0] meta_table_io_data_in_a_field_type_30_sub_class_id; // @[XRam.scala 102:23]
  wire  meta_table_io_data_in_a_field_type_30_is_host; // @[XRam.scala 102:23]
  wire  meta_table_io_data_in_a_field_type_31_is_repeated; // @[XRam.scala 102:23]
  wire [4:0] meta_table_io_data_in_a_field_type_31_field_type; // @[XRam.scala 102:23]
  wire [15:0] meta_table_io_data_in_a_field_type_31_sub_class_id; // @[XRam.scala 102:23]
  wire  meta_table_io_data_in_a_field_type_31_is_host; // @[XRam.scala 102:23]
  wire  meta_table_io_data_in_a_field_type_32_is_repeated; // @[XRam.scala 102:23]
  wire [4:0] meta_table_io_data_in_a_field_type_32_field_type; // @[XRam.scala 102:23]
  wire [15:0] meta_table_io_data_in_a_field_type_32_sub_class_id; // @[XRam.scala 102:23]
  wire  meta_table_io_data_in_a_field_type_32_is_host; // @[XRam.scala 102:23]
  wire [7:0] meta_table_io_data_out_b_max_field_num; // @[XRam.scala 102:23]
  wire  meta_table_io_data_out_b_field_type_0_is_repeated; // @[XRam.scala 102:23]
  wire [4:0] meta_table_io_data_out_b_field_type_0_field_type; // @[XRam.scala 102:23]
  wire [15:0] meta_table_io_data_out_b_field_type_0_sub_class_id; // @[XRam.scala 102:23]
  wire  meta_table_io_data_out_b_field_type_1_is_repeated; // @[XRam.scala 102:23]
  wire [4:0] meta_table_io_data_out_b_field_type_1_field_type; // @[XRam.scala 102:23]
  wire [15:0] meta_table_io_data_out_b_field_type_1_sub_class_id; // @[XRam.scala 102:23]
  wire  meta_table_io_data_out_b_field_type_2_is_repeated; // @[XRam.scala 102:23]
  wire [4:0] meta_table_io_data_out_b_field_type_2_field_type; // @[XRam.scala 102:23]
  wire [15:0] meta_table_io_data_out_b_field_type_2_sub_class_id; // @[XRam.scala 102:23]
  wire  meta_table_io_data_out_b_field_type_3_is_repeated; // @[XRam.scala 102:23]
  wire [4:0] meta_table_io_data_out_b_field_type_3_field_type; // @[XRam.scala 102:23]
  wire [15:0] meta_table_io_data_out_b_field_type_3_sub_class_id; // @[XRam.scala 102:23]
  wire  meta_table_io_data_out_b_field_type_4_is_repeated; // @[XRam.scala 102:23]
  wire [4:0] meta_table_io_data_out_b_field_type_4_field_type; // @[XRam.scala 102:23]
  wire [15:0] meta_table_io_data_out_b_field_type_4_sub_class_id; // @[XRam.scala 102:23]
  wire  meta_table_io_data_out_b_field_type_5_is_repeated; // @[XRam.scala 102:23]
  wire [4:0] meta_table_io_data_out_b_field_type_5_field_type; // @[XRam.scala 102:23]
  wire [15:0] meta_table_io_data_out_b_field_type_5_sub_class_id; // @[XRam.scala 102:23]
  wire  meta_table_io_data_out_b_field_type_6_is_repeated; // @[XRam.scala 102:23]
  wire [4:0] meta_table_io_data_out_b_field_type_6_field_type; // @[XRam.scala 102:23]
  wire [15:0] meta_table_io_data_out_b_field_type_6_sub_class_id; // @[XRam.scala 102:23]
  wire  meta_table_io_data_out_b_field_type_7_is_repeated; // @[XRam.scala 102:23]
  wire [4:0] meta_table_io_data_out_b_field_type_7_field_type; // @[XRam.scala 102:23]
  wire [15:0] meta_table_io_data_out_b_field_type_7_sub_class_id; // @[XRam.scala 102:23]
  wire  meta_table_io_data_out_b_field_type_8_is_repeated; // @[XRam.scala 102:23]
  wire [4:0] meta_table_io_data_out_b_field_type_8_field_type; // @[XRam.scala 102:23]
  wire [15:0] meta_table_io_data_out_b_field_type_8_sub_class_id; // @[XRam.scala 102:23]
  wire  meta_table_io_data_out_b_field_type_9_is_repeated; // @[XRam.scala 102:23]
  wire [4:0] meta_table_io_data_out_b_field_type_9_field_type; // @[XRam.scala 102:23]
  wire [15:0] meta_table_io_data_out_b_field_type_9_sub_class_id; // @[XRam.scala 102:23]
  wire  meta_table_io_data_out_b_field_type_10_is_repeated; // @[XRam.scala 102:23]
  wire [4:0] meta_table_io_data_out_b_field_type_10_field_type; // @[XRam.scala 102:23]
  wire [15:0] meta_table_io_data_out_b_field_type_10_sub_class_id; // @[XRam.scala 102:23]
  wire  meta_table_io_data_out_b_field_type_11_is_repeated; // @[XRam.scala 102:23]
  wire [4:0] meta_table_io_data_out_b_field_type_11_field_type; // @[XRam.scala 102:23]
  wire [15:0] meta_table_io_data_out_b_field_type_11_sub_class_id; // @[XRam.scala 102:23]
  wire  meta_table_io_data_out_b_field_type_12_is_repeated; // @[XRam.scala 102:23]
  wire [4:0] meta_table_io_data_out_b_field_type_12_field_type; // @[XRam.scala 102:23]
  wire [15:0] meta_table_io_data_out_b_field_type_12_sub_class_id; // @[XRam.scala 102:23]
  wire  meta_table_io_data_out_b_field_type_13_is_repeated; // @[XRam.scala 102:23]
  wire [4:0] meta_table_io_data_out_b_field_type_13_field_type; // @[XRam.scala 102:23]
  wire [15:0] meta_table_io_data_out_b_field_type_13_sub_class_id; // @[XRam.scala 102:23]
  wire  meta_table_io_data_out_b_field_type_14_is_repeated; // @[XRam.scala 102:23]
  wire [4:0] meta_table_io_data_out_b_field_type_14_field_type; // @[XRam.scala 102:23]
  wire [15:0] meta_table_io_data_out_b_field_type_14_sub_class_id; // @[XRam.scala 102:23]
  wire  meta_table_io_data_out_b_field_type_15_is_repeated; // @[XRam.scala 102:23]
  wire [4:0] meta_table_io_data_out_b_field_type_15_field_type; // @[XRam.scala 102:23]
  wire [15:0] meta_table_io_data_out_b_field_type_15_sub_class_id; // @[XRam.scala 102:23]
  wire  meta_table_io_data_out_b_field_type_16_is_repeated; // @[XRam.scala 102:23]
  wire [4:0] meta_table_io_data_out_b_field_type_16_field_type; // @[XRam.scala 102:23]
  wire [15:0] meta_table_io_data_out_b_field_type_16_sub_class_id; // @[XRam.scala 102:23]
  wire  meta_table_io_data_out_b_field_type_17_is_repeated; // @[XRam.scala 102:23]
  wire [4:0] meta_table_io_data_out_b_field_type_17_field_type; // @[XRam.scala 102:23]
  wire [15:0] meta_table_io_data_out_b_field_type_17_sub_class_id; // @[XRam.scala 102:23]
  wire  meta_table_io_data_out_b_field_type_18_is_repeated; // @[XRam.scala 102:23]
  wire [4:0] meta_table_io_data_out_b_field_type_18_field_type; // @[XRam.scala 102:23]
  wire [15:0] meta_table_io_data_out_b_field_type_18_sub_class_id; // @[XRam.scala 102:23]
  wire  meta_table_io_data_out_b_field_type_19_is_repeated; // @[XRam.scala 102:23]
  wire [4:0] meta_table_io_data_out_b_field_type_19_field_type; // @[XRam.scala 102:23]
  wire [15:0] meta_table_io_data_out_b_field_type_19_sub_class_id; // @[XRam.scala 102:23]
  wire  meta_table_io_data_out_b_field_type_20_is_repeated; // @[XRam.scala 102:23]
  wire [4:0] meta_table_io_data_out_b_field_type_20_field_type; // @[XRam.scala 102:23]
  wire [15:0] meta_table_io_data_out_b_field_type_20_sub_class_id; // @[XRam.scala 102:23]
  wire  meta_table_io_data_out_b_field_type_21_is_repeated; // @[XRam.scala 102:23]
  wire [4:0] meta_table_io_data_out_b_field_type_21_field_type; // @[XRam.scala 102:23]
  wire [15:0] meta_table_io_data_out_b_field_type_21_sub_class_id; // @[XRam.scala 102:23]
  wire  meta_table_io_data_out_b_field_type_22_is_repeated; // @[XRam.scala 102:23]
  wire [4:0] meta_table_io_data_out_b_field_type_22_field_type; // @[XRam.scala 102:23]
  wire [15:0] meta_table_io_data_out_b_field_type_22_sub_class_id; // @[XRam.scala 102:23]
  wire  meta_table_io_data_out_b_field_type_23_is_repeated; // @[XRam.scala 102:23]
  wire [4:0] meta_table_io_data_out_b_field_type_23_field_type; // @[XRam.scala 102:23]
  wire [15:0] meta_table_io_data_out_b_field_type_23_sub_class_id; // @[XRam.scala 102:23]
  wire  meta_table_io_data_out_b_field_type_24_is_repeated; // @[XRam.scala 102:23]
  wire [4:0] meta_table_io_data_out_b_field_type_24_field_type; // @[XRam.scala 102:23]
  wire [15:0] meta_table_io_data_out_b_field_type_24_sub_class_id; // @[XRam.scala 102:23]
  wire  meta_table_io_data_out_b_field_type_25_is_repeated; // @[XRam.scala 102:23]
  wire [4:0] meta_table_io_data_out_b_field_type_25_field_type; // @[XRam.scala 102:23]
  wire [15:0] meta_table_io_data_out_b_field_type_25_sub_class_id; // @[XRam.scala 102:23]
  wire  meta_table_io_data_out_b_field_type_26_is_repeated; // @[XRam.scala 102:23]
  wire [4:0] meta_table_io_data_out_b_field_type_26_field_type; // @[XRam.scala 102:23]
  wire [15:0] meta_table_io_data_out_b_field_type_26_sub_class_id; // @[XRam.scala 102:23]
  wire  meta_table_io_data_out_b_field_type_27_is_repeated; // @[XRam.scala 102:23]
  wire [4:0] meta_table_io_data_out_b_field_type_27_field_type; // @[XRam.scala 102:23]
  wire [15:0] meta_table_io_data_out_b_field_type_27_sub_class_id; // @[XRam.scala 102:23]
  wire  meta_table_io_data_out_b_field_type_28_is_repeated; // @[XRam.scala 102:23]
  wire [4:0] meta_table_io_data_out_b_field_type_28_field_type; // @[XRam.scala 102:23]
  wire [15:0] meta_table_io_data_out_b_field_type_28_sub_class_id; // @[XRam.scala 102:23]
  wire  meta_table_io_data_out_b_field_type_29_is_repeated; // @[XRam.scala 102:23]
  wire [4:0] meta_table_io_data_out_b_field_type_29_field_type; // @[XRam.scala 102:23]
  wire [15:0] meta_table_io_data_out_b_field_type_29_sub_class_id; // @[XRam.scala 102:23]
  wire  meta_table_io_data_out_b_field_type_30_is_repeated; // @[XRam.scala 102:23]
  wire [4:0] meta_table_io_data_out_b_field_type_30_field_type; // @[XRam.scala 102:23]
  wire [15:0] meta_table_io_data_out_b_field_type_30_sub_class_id; // @[XRam.scala 102:23]
  wire  meta_table_io_data_out_b_field_type_31_is_repeated; // @[XRam.scala 102:23]
  wire [4:0] meta_table_io_data_out_b_field_type_31_field_type; // @[XRam.scala 102:23]
  wire [15:0] meta_table_io_data_out_b_field_type_31_sub_class_id; // @[XRam.scala 102:23]
  wire  meta_table_io_data_out_b_field_type_32_is_repeated; // @[XRam.scala 102:23]
  wire [4:0] meta_table_io_data_out_b_field_type_32_field_type; // @[XRam.scala 102:23]
  wire [15:0] meta_table_io_data_out_b_field_type_32_sub_class_id; // @[XRam.scala 102:23]
  reg [31:0] counter; // @[Collector.scala 169:42]
  wire  _T = io_class_meta_init_ready & io_class_meta_init_valid; // @[Decoupled.scala 40:37]
  wire [31:0] _counter_T_1 = counter + 32'h1; // @[Collector.scala 171:51]
  reg [1:0] state; // @[ClassMetaTable.scala 67:46]
  wire  _s_class_meta_req_fifo_io_out_ready_T_1 = ~io_class_meta_init_valid; // @[ClassMetaTable.scala 74:54]
  wire  _s_class_meta_req_fifo_io_out_ready_T_2 = state == 2'h0; // @[ClassMetaTable.scala 74:97]
  wire  _T_2 = s_class_meta_req_fifo_io_out_ready & s_class_meta_req_fifo_io_out_valid; // @[Decoupled.scala 40:37]
  wire  _T_3 = d_class_meta_req_fifo_io_out_ready & d_class_meta_req_fifo_io_out_valid; // @[Decoupled.scala 40:37]
  wire [9:0] _GEN_1 = _T_3 ? d_class_meta_req_fifo_io_out_bits_class_id : 10'h0; // @[ClassMetaTable.scala 94:52 ClassMetaTable.scala 95:49 ClassMetaTable.scala 70:42]
  wire [9:0] _GEN_4 = _T_2 ? s_class_meta_req_fifo_io_out_bits_class_id : _GEN_1; // @[ClassMetaTable.scala 90:52 ClassMetaTable.scala 91:49]
  XQueue_4 s_class_meta_req_fifo ( // @[XQueue.scala 35:23]
    .clock(s_class_meta_req_fifo_clock),
    .reset(s_class_meta_req_fifo_reset),
    .io_in_ready(s_class_meta_req_fifo_io_in_ready),
    .io_in_valid(s_class_meta_req_fifo_io_in_valid),
    .io_in_bits_class_id(s_class_meta_req_fifo_io_in_bits_class_id),
    .io_out_ready(s_class_meta_req_fifo_io_out_ready),
    .io_out_valid(s_class_meta_req_fifo_io_out_valid),
    .io_out_bits_class_id(s_class_meta_req_fifo_io_out_bits_class_id)
  );
  XQueue_4 d_class_meta_req_fifo ( // @[XQueue.scala 35:23]
    .clock(d_class_meta_req_fifo_clock),
    .reset(d_class_meta_req_fifo_reset),
    .io_in_ready(d_class_meta_req_fifo_io_in_ready),
    .io_in_valid(d_class_meta_req_fifo_io_in_valid),
    .io_in_bits_class_id(d_class_meta_req_fifo_io_in_bits_class_id),
    .io_out_ready(d_class_meta_req_fifo_io_out_ready),
    .io_out_valid(d_class_meta_req_fifo_io_out_valid),
    .io_out_bits_class_id(d_class_meta_req_fifo_io_out_bits_class_id)
  );
  XRam_1 meta_table ( // @[XRam.scala 102:23]
    .clock(meta_table_clock),
    .reset(meta_table_reset),
    .io_addr_a(meta_table_io_addr_a),
    .io_addr_b(meta_table_io_addr_b),
    .io_wr_en_a(meta_table_io_wr_en_a),
    .io_data_in_a_class_length(meta_table_io_data_in_a_class_length),
    .io_data_in_a_max_field_num(meta_table_io_data_in_a_max_field_num),
    .io_data_in_a_field_type_0_is_repeated(meta_table_io_data_in_a_field_type_0_is_repeated),
    .io_data_in_a_field_type_0_field_type(meta_table_io_data_in_a_field_type_0_field_type),
    .io_data_in_a_field_type_0_sub_class_id(meta_table_io_data_in_a_field_type_0_sub_class_id),
    .io_data_in_a_field_type_0_is_host(meta_table_io_data_in_a_field_type_0_is_host),
    .io_data_in_a_field_type_1_is_repeated(meta_table_io_data_in_a_field_type_1_is_repeated),
    .io_data_in_a_field_type_1_field_type(meta_table_io_data_in_a_field_type_1_field_type),
    .io_data_in_a_field_type_1_sub_class_id(meta_table_io_data_in_a_field_type_1_sub_class_id),
    .io_data_in_a_field_type_1_is_host(meta_table_io_data_in_a_field_type_1_is_host),
    .io_data_in_a_field_type_2_is_repeated(meta_table_io_data_in_a_field_type_2_is_repeated),
    .io_data_in_a_field_type_2_field_type(meta_table_io_data_in_a_field_type_2_field_type),
    .io_data_in_a_field_type_2_sub_class_id(meta_table_io_data_in_a_field_type_2_sub_class_id),
    .io_data_in_a_field_type_2_is_host(meta_table_io_data_in_a_field_type_2_is_host),
    .io_data_in_a_field_type_3_is_repeated(meta_table_io_data_in_a_field_type_3_is_repeated),
    .io_data_in_a_field_type_3_field_type(meta_table_io_data_in_a_field_type_3_field_type),
    .io_data_in_a_field_type_3_sub_class_id(meta_table_io_data_in_a_field_type_3_sub_class_id),
    .io_data_in_a_field_type_3_is_host(meta_table_io_data_in_a_field_type_3_is_host),
    .io_data_in_a_field_type_4_is_repeated(meta_table_io_data_in_a_field_type_4_is_repeated),
    .io_data_in_a_field_type_4_field_type(meta_table_io_data_in_a_field_type_4_field_type),
    .io_data_in_a_field_type_4_sub_class_id(meta_table_io_data_in_a_field_type_4_sub_class_id),
    .io_data_in_a_field_type_4_is_host(meta_table_io_data_in_a_field_type_4_is_host),
    .io_data_in_a_field_type_5_is_repeated(meta_table_io_data_in_a_field_type_5_is_repeated),
    .io_data_in_a_field_type_5_field_type(meta_table_io_data_in_a_field_type_5_field_type),
    .io_data_in_a_field_type_5_sub_class_id(meta_table_io_data_in_a_field_type_5_sub_class_id),
    .io_data_in_a_field_type_5_is_host(meta_table_io_data_in_a_field_type_5_is_host),
    .io_data_in_a_field_type_6_is_repeated(meta_table_io_data_in_a_field_type_6_is_repeated),
    .io_data_in_a_field_type_6_field_type(meta_table_io_data_in_a_field_type_6_field_type),
    .io_data_in_a_field_type_6_sub_class_id(meta_table_io_data_in_a_field_type_6_sub_class_id),
    .io_data_in_a_field_type_6_is_host(meta_table_io_data_in_a_field_type_6_is_host),
    .io_data_in_a_field_type_7_is_repeated(meta_table_io_data_in_a_field_type_7_is_repeated),
    .io_data_in_a_field_type_7_field_type(meta_table_io_data_in_a_field_type_7_field_type),
    .io_data_in_a_field_type_7_sub_class_id(meta_table_io_data_in_a_field_type_7_sub_class_id),
    .io_data_in_a_field_type_7_is_host(meta_table_io_data_in_a_field_type_7_is_host),
    .io_data_in_a_field_type_8_is_repeated(meta_table_io_data_in_a_field_type_8_is_repeated),
    .io_data_in_a_field_type_8_field_type(meta_table_io_data_in_a_field_type_8_field_type),
    .io_data_in_a_field_type_8_sub_class_id(meta_table_io_data_in_a_field_type_8_sub_class_id),
    .io_data_in_a_field_type_8_is_host(meta_table_io_data_in_a_field_type_8_is_host),
    .io_data_in_a_field_type_9_is_repeated(meta_table_io_data_in_a_field_type_9_is_repeated),
    .io_data_in_a_field_type_9_field_type(meta_table_io_data_in_a_field_type_9_field_type),
    .io_data_in_a_field_type_9_sub_class_id(meta_table_io_data_in_a_field_type_9_sub_class_id),
    .io_data_in_a_field_type_9_is_host(meta_table_io_data_in_a_field_type_9_is_host),
    .io_data_in_a_field_type_10_is_repeated(meta_table_io_data_in_a_field_type_10_is_repeated),
    .io_data_in_a_field_type_10_field_type(meta_table_io_data_in_a_field_type_10_field_type),
    .io_data_in_a_field_type_10_sub_class_id(meta_table_io_data_in_a_field_type_10_sub_class_id),
    .io_data_in_a_field_type_10_is_host(meta_table_io_data_in_a_field_type_10_is_host),
    .io_data_in_a_field_type_11_is_repeated(meta_table_io_data_in_a_field_type_11_is_repeated),
    .io_data_in_a_field_type_11_field_type(meta_table_io_data_in_a_field_type_11_field_type),
    .io_data_in_a_field_type_11_sub_class_id(meta_table_io_data_in_a_field_type_11_sub_class_id),
    .io_data_in_a_field_type_11_is_host(meta_table_io_data_in_a_field_type_11_is_host),
    .io_data_in_a_field_type_12_is_repeated(meta_table_io_data_in_a_field_type_12_is_repeated),
    .io_data_in_a_field_type_12_field_type(meta_table_io_data_in_a_field_type_12_field_type),
    .io_data_in_a_field_type_12_sub_class_id(meta_table_io_data_in_a_field_type_12_sub_class_id),
    .io_data_in_a_field_type_12_is_host(meta_table_io_data_in_a_field_type_12_is_host),
    .io_data_in_a_field_type_13_is_repeated(meta_table_io_data_in_a_field_type_13_is_repeated),
    .io_data_in_a_field_type_13_field_type(meta_table_io_data_in_a_field_type_13_field_type),
    .io_data_in_a_field_type_13_sub_class_id(meta_table_io_data_in_a_field_type_13_sub_class_id),
    .io_data_in_a_field_type_13_is_host(meta_table_io_data_in_a_field_type_13_is_host),
    .io_data_in_a_field_type_14_is_repeated(meta_table_io_data_in_a_field_type_14_is_repeated),
    .io_data_in_a_field_type_14_field_type(meta_table_io_data_in_a_field_type_14_field_type),
    .io_data_in_a_field_type_14_sub_class_id(meta_table_io_data_in_a_field_type_14_sub_class_id),
    .io_data_in_a_field_type_14_is_host(meta_table_io_data_in_a_field_type_14_is_host),
    .io_data_in_a_field_type_15_is_repeated(meta_table_io_data_in_a_field_type_15_is_repeated),
    .io_data_in_a_field_type_15_field_type(meta_table_io_data_in_a_field_type_15_field_type),
    .io_data_in_a_field_type_15_sub_class_id(meta_table_io_data_in_a_field_type_15_sub_class_id),
    .io_data_in_a_field_type_15_is_host(meta_table_io_data_in_a_field_type_15_is_host),
    .io_data_in_a_field_type_16_is_repeated(meta_table_io_data_in_a_field_type_16_is_repeated),
    .io_data_in_a_field_type_16_field_type(meta_table_io_data_in_a_field_type_16_field_type),
    .io_data_in_a_field_type_16_sub_class_id(meta_table_io_data_in_a_field_type_16_sub_class_id),
    .io_data_in_a_field_type_16_is_host(meta_table_io_data_in_a_field_type_16_is_host),
    .io_data_in_a_field_type_17_is_repeated(meta_table_io_data_in_a_field_type_17_is_repeated),
    .io_data_in_a_field_type_17_field_type(meta_table_io_data_in_a_field_type_17_field_type),
    .io_data_in_a_field_type_17_sub_class_id(meta_table_io_data_in_a_field_type_17_sub_class_id),
    .io_data_in_a_field_type_17_is_host(meta_table_io_data_in_a_field_type_17_is_host),
    .io_data_in_a_field_type_18_is_repeated(meta_table_io_data_in_a_field_type_18_is_repeated),
    .io_data_in_a_field_type_18_field_type(meta_table_io_data_in_a_field_type_18_field_type),
    .io_data_in_a_field_type_18_sub_class_id(meta_table_io_data_in_a_field_type_18_sub_class_id),
    .io_data_in_a_field_type_18_is_host(meta_table_io_data_in_a_field_type_18_is_host),
    .io_data_in_a_field_type_19_is_repeated(meta_table_io_data_in_a_field_type_19_is_repeated),
    .io_data_in_a_field_type_19_field_type(meta_table_io_data_in_a_field_type_19_field_type),
    .io_data_in_a_field_type_19_sub_class_id(meta_table_io_data_in_a_field_type_19_sub_class_id),
    .io_data_in_a_field_type_19_is_host(meta_table_io_data_in_a_field_type_19_is_host),
    .io_data_in_a_field_type_20_is_repeated(meta_table_io_data_in_a_field_type_20_is_repeated),
    .io_data_in_a_field_type_20_field_type(meta_table_io_data_in_a_field_type_20_field_type),
    .io_data_in_a_field_type_20_sub_class_id(meta_table_io_data_in_a_field_type_20_sub_class_id),
    .io_data_in_a_field_type_20_is_host(meta_table_io_data_in_a_field_type_20_is_host),
    .io_data_in_a_field_type_21_is_repeated(meta_table_io_data_in_a_field_type_21_is_repeated),
    .io_data_in_a_field_type_21_field_type(meta_table_io_data_in_a_field_type_21_field_type),
    .io_data_in_a_field_type_21_sub_class_id(meta_table_io_data_in_a_field_type_21_sub_class_id),
    .io_data_in_a_field_type_21_is_host(meta_table_io_data_in_a_field_type_21_is_host),
    .io_data_in_a_field_type_22_is_repeated(meta_table_io_data_in_a_field_type_22_is_repeated),
    .io_data_in_a_field_type_22_field_type(meta_table_io_data_in_a_field_type_22_field_type),
    .io_data_in_a_field_type_22_sub_class_id(meta_table_io_data_in_a_field_type_22_sub_class_id),
    .io_data_in_a_field_type_22_is_host(meta_table_io_data_in_a_field_type_22_is_host),
    .io_data_in_a_field_type_23_is_repeated(meta_table_io_data_in_a_field_type_23_is_repeated),
    .io_data_in_a_field_type_23_field_type(meta_table_io_data_in_a_field_type_23_field_type),
    .io_data_in_a_field_type_23_sub_class_id(meta_table_io_data_in_a_field_type_23_sub_class_id),
    .io_data_in_a_field_type_23_is_host(meta_table_io_data_in_a_field_type_23_is_host),
    .io_data_in_a_field_type_24_is_repeated(meta_table_io_data_in_a_field_type_24_is_repeated),
    .io_data_in_a_field_type_24_field_type(meta_table_io_data_in_a_field_type_24_field_type),
    .io_data_in_a_field_type_24_sub_class_id(meta_table_io_data_in_a_field_type_24_sub_class_id),
    .io_data_in_a_field_type_24_is_host(meta_table_io_data_in_a_field_type_24_is_host),
    .io_data_in_a_field_type_25_is_repeated(meta_table_io_data_in_a_field_type_25_is_repeated),
    .io_data_in_a_field_type_25_field_type(meta_table_io_data_in_a_field_type_25_field_type),
    .io_data_in_a_field_type_25_sub_class_id(meta_table_io_data_in_a_field_type_25_sub_class_id),
    .io_data_in_a_field_type_25_is_host(meta_table_io_data_in_a_field_type_25_is_host),
    .io_data_in_a_field_type_26_is_repeated(meta_table_io_data_in_a_field_type_26_is_repeated),
    .io_data_in_a_field_type_26_field_type(meta_table_io_data_in_a_field_type_26_field_type),
    .io_data_in_a_field_type_26_sub_class_id(meta_table_io_data_in_a_field_type_26_sub_class_id),
    .io_data_in_a_field_type_26_is_host(meta_table_io_data_in_a_field_type_26_is_host),
    .io_data_in_a_field_type_27_is_repeated(meta_table_io_data_in_a_field_type_27_is_repeated),
    .io_data_in_a_field_type_27_field_type(meta_table_io_data_in_a_field_type_27_field_type),
    .io_data_in_a_field_type_27_sub_class_id(meta_table_io_data_in_a_field_type_27_sub_class_id),
    .io_data_in_a_field_type_27_is_host(meta_table_io_data_in_a_field_type_27_is_host),
    .io_data_in_a_field_type_28_is_repeated(meta_table_io_data_in_a_field_type_28_is_repeated),
    .io_data_in_a_field_type_28_field_type(meta_table_io_data_in_a_field_type_28_field_type),
    .io_data_in_a_field_type_28_sub_class_id(meta_table_io_data_in_a_field_type_28_sub_class_id),
    .io_data_in_a_field_type_28_is_host(meta_table_io_data_in_a_field_type_28_is_host),
    .io_data_in_a_field_type_29_is_repeated(meta_table_io_data_in_a_field_type_29_is_repeated),
    .io_data_in_a_field_type_29_field_type(meta_table_io_data_in_a_field_type_29_field_type),
    .io_data_in_a_field_type_29_sub_class_id(meta_table_io_data_in_a_field_type_29_sub_class_id),
    .io_data_in_a_field_type_29_is_host(meta_table_io_data_in_a_field_type_29_is_host),
    .io_data_in_a_field_type_30_is_repeated(meta_table_io_data_in_a_field_type_30_is_repeated),
    .io_data_in_a_field_type_30_field_type(meta_table_io_data_in_a_field_type_30_field_type),
    .io_data_in_a_field_type_30_sub_class_id(meta_table_io_data_in_a_field_type_30_sub_class_id),
    .io_data_in_a_field_type_30_is_host(meta_table_io_data_in_a_field_type_30_is_host),
    .io_data_in_a_field_type_31_is_repeated(meta_table_io_data_in_a_field_type_31_is_repeated),
    .io_data_in_a_field_type_31_field_type(meta_table_io_data_in_a_field_type_31_field_type),
    .io_data_in_a_field_type_31_sub_class_id(meta_table_io_data_in_a_field_type_31_sub_class_id),
    .io_data_in_a_field_type_31_is_host(meta_table_io_data_in_a_field_type_31_is_host),
    .io_data_in_a_field_type_32_is_repeated(meta_table_io_data_in_a_field_type_32_is_repeated),
    .io_data_in_a_field_type_32_field_type(meta_table_io_data_in_a_field_type_32_field_type),
    .io_data_in_a_field_type_32_sub_class_id(meta_table_io_data_in_a_field_type_32_sub_class_id),
    .io_data_in_a_field_type_32_is_host(meta_table_io_data_in_a_field_type_32_is_host),
    .io_data_out_b_max_field_num(meta_table_io_data_out_b_max_field_num),
    .io_data_out_b_field_type_0_is_repeated(meta_table_io_data_out_b_field_type_0_is_repeated),
    .io_data_out_b_field_type_0_field_type(meta_table_io_data_out_b_field_type_0_field_type),
    .io_data_out_b_field_type_0_sub_class_id(meta_table_io_data_out_b_field_type_0_sub_class_id),
    .io_data_out_b_field_type_1_is_repeated(meta_table_io_data_out_b_field_type_1_is_repeated),
    .io_data_out_b_field_type_1_field_type(meta_table_io_data_out_b_field_type_1_field_type),
    .io_data_out_b_field_type_1_sub_class_id(meta_table_io_data_out_b_field_type_1_sub_class_id),
    .io_data_out_b_field_type_2_is_repeated(meta_table_io_data_out_b_field_type_2_is_repeated),
    .io_data_out_b_field_type_2_field_type(meta_table_io_data_out_b_field_type_2_field_type),
    .io_data_out_b_field_type_2_sub_class_id(meta_table_io_data_out_b_field_type_2_sub_class_id),
    .io_data_out_b_field_type_3_is_repeated(meta_table_io_data_out_b_field_type_3_is_repeated),
    .io_data_out_b_field_type_3_field_type(meta_table_io_data_out_b_field_type_3_field_type),
    .io_data_out_b_field_type_3_sub_class_id(meta_table_io_data_out_b_field_type_3_sub_class_id),
    .io_data_out_b_field_type_4_is_repeated(meta_table_io_data_out_b_field_type_4_is_repeated),
    .io_data_out_b_field_type_4_field_type(meta_table_io_data_out_b_field_type_4_field_type),
    .io_data_out_b_field_type_4_sub_class_id(meta_table_io_data_out_b_field_type_4_sub_class_id),
    .io_data_out_b_field_type_5_is_repeated(meta_table_io_data_out_b_field_type_5_is_repeated),
    .io_data_out_b_field_type_5_field_type(meta_table_io_data_out_b_field_type_5_field_type),
    .io_data_out_b_field_type_5_sub_class_id(meta_table_io_data_out_b_field_type_5_sub_class_id),
    .io_data_out_b_field_type_6_is_repeated(meta_table_io_data_out_b_field_type_6_is_repeated),
    .io_data_out_b_field_type_6_field_type(meta_table_io_data_out_b_field_type_6_field_type),
    .io_data_out_b_field_type_6_sub_class_id(meta_table_io_data_out_b_field_type_6_sub_class_id),
    .io_data_out_b_field_type_7_is_repeated(meta_table_io_data_out_b_field_type_7_is_repeated),
    .io_data_out_b_field_type_7_field_type(meta_table_io_data_out_b_field_type_7_field_type),
    .io_data_out_b_field_type_7_sub_class_id(meta_table_io_data_out_b_field_type_7_sub_class_id),
    .io_data_out_b_field_type_8_is_repeated(meta_table_io_data_out_b_field_type_8_is_repeated),
    .io_data_out_b_field_type_8_field_type(meta_table_io_data_out_b_field_type_8_field_type),
    .io_data_out_b_field_type_8_sub_class_id(meta_table_io_data_out_b_field_type_8_sub_class_id),
    .io_data_out_b_field_type_9_is_repeated(meta_table_io_data_out_b_field_type_9_is_repeated),
    .io_data_out_b_field_type_9_field_type(meta_table_io_data_out_b_field_type_9_field_type),
    .io_data_out_b_field_type_9_sub_class_id(meta_table_io_data_out_b_field_type_9_sub_class_id),
    .io_data_out_b_field_type_10_is_repeated(meta_table_io_data_out_b_field_type_10_is_repeated),
    .io_data_out_b_field_type_10_field_type(meta_table_io_data_out_b_field_type_10_field_type),
    .io_data_out_b_field_type_10_sub_class_id(meta_table_io_data_out_b_field_type_10_sub_class_id),
    .io_data_out_b_field_type_11_is_repeated(meta_table_io_data_out_b_field_type_11_is_repeated),
    .io_data_out_b_field_type_11_field_type(meta_table_io_data_out_b_field_type_11_field_type),
    .io_data_out_b_field_type_11_sub_class_id(meta_table_io_data_out_b_field_type_11_sub_class_id),
    .io_data_out_b_field_type_12_is_repeated(meta_table_io_data_out_b_field_type_12_is_repeated),
    .io_data_out_b_field_type_12_field_type(meta_table_io_data_out_b_field_type_12_field_type),
    .io_data_out_b_field_type_12_sub_class_id(meta_table_io_data_out_b_field_type_12_sub_class_id),
    .io_data_out_b_field_type_13_is_repeated(meta_table_io_data_out_b_field_type_13_is_repeated),
    .io_data_out_b_field_type_13_field_type(meta_table_io_data_out_b_field_type_13_field_type),
    .io_data_out_b_field_type_13_sub_class_id(meta_table_io_data_out_b_field_type_13_sub_class_id),
    .io_data_out_b_field_type_14_is_repeated(meta_table_io_data_out_b_field_type_14_is_repeated),
    .io_data_out_b_field_type_14_field_type(meta_table_io_data_out_b_field_type_14_field_type),
    .io_data_out_b_field_type_14_sub_class_id(meta_table_io_data_out_b_field_type_14_sub_class_id),
    .io_data_out_b_field_type_15_is_repeated(meta_table_io_data_out_b_field_type_15_is_repeated),
    .io_data_out_b_field_type_15_field_type(meta_table_io_data_out_b_field_type_15_field_type),
    .io_data_out_b_field_type_15_sub_class_id(meta_table_io_data_out_b_field_type_15_sub_class_id),
    .io_data_out_b_field_type_16_is_repeated(meta_table_io_data_out_b_field_type_16_is_repeated),
    .io_data_out_b_field_type_16_field_type(meta_table_io_data_out_b_field_type_16_field_type),
    .io_data_out_b_field_type_16_sub_class_id(meta_table_io_data_out_b_field_type_16_sub_class_id),
    .io_data_out_b_field_type_17_is_repeated(meta_table_io_data_out_b_field_type_17_is_repeated),
    .io_data_out_b_field_type_17_field_type(meta_table_io_data_out_b_field_type_17_field_type),
    .io_data_out_b_field_type_17_sub_class_id(meta_table_io_data_out_b_field_type_17_sub_class_id),
    .io_data_out_b_field_type_18_is_repeated(meta_table_io_data_out_b_field_type_18_is_repeated),
    .io_data_out_b_field_type_18_field_type(meta_table_io_data_out_b_field_type_18_field_type),
    .io_data_out_b_field_type_18_sub_class_id(meta_table_io_data_out_b_field_type_18_sub_class_id),
    .io_data_out_b_field_type_19_is_repeated(meta_table_io_data_out_b_field_type_19_is_repeated),
    .io_data_out_b_field_type_19_field_type(meta_table_io_data_out_b_field_type_19_field_type),
    .io_data_out_b_field_type_19_sub_class_id(meta_table_io_data_out_b_field_type_19_sub_class_id),
    .io_data_out_b_field_type_20_is_repeated(meta_table_io_data_out_b_field_type_20_is_repeated),
    .io_data_out_b_field_type_20_field_type(meta_table_io_data_out_b_field_type_20_field_type),
    .io_data_out_b_field_type_20_sub_class_id(meta_table_io_data_out_b_field_type_20_sub_class_id),
    .io_data_out_b_field_type_21_is_repeated(meta_table_io_data_out_b_field_type_21_is_repeated),
    .io_data_out_b_field_type_21_field_type(meta_table_io_data_out_b_field_type_21_field_type),
    .io_data_out_b_field_type_21_sub_class_id(meta_table_io_data_out_b_field_type_21_sub_class_id),
    .io_data_out_b_field_type_22_is_repeated(meta_table_io_data_out_b_field_type_22_is_repeated),
    .io_data_out_b_field_type_22_field_type(meta_table_io_data_out_b_field_type_22_field_type),
    .io_data_out_b_field_type_22_sub_class_id(meta_table_io_data_out_b_field_type_22_sub_class_id),
    .io_data_out_b_field_type_23_is_repeated(meta_table_io_data_out_b_field_type_23_is_repeated),
    .io_data_out_b_field_type_23_field_type(meta_table_io_data_out_b_field_type_23_field_type),
    .io_data_out_b_field_type_23_sub_class_id(meta_table_io_data_out_b_field_type_23_sub_class_id),
    .io_data_out_b_field_type_24_is_repeated(meta_table_io_data_out_b_field_type_24_is_repeated),
    .io_data_out_b_field_type_24_field_type(meta_table_io_data_out_b_field_type_24_field_type),
    .io_data_out_b_field_type_24_sub_class_id(meta_table_io_data_out_b_field_type_24_sub_class_id),
    .io_data_out_b_field_type_25_is_repeated(meta_table_io_data_out_b_field_type_25_is_repeated),
    .io_data_out_b_field_type_25_field_type(meta_table_io_data_out_b_field_type_25_field_type),
    .io_data_out_b_field_type_25_sub_class_id(meta_table_io_data_out_b_field_type_25_sub_class_id),
    .io_data_out_b_field_type_26_is_repeated(meta_table_io_data_out_b_field_type_26_is_repeated),
    .io_data_out_b_field_type_26_field_type(meta_table_io_data_out_b_field_type_26_field_type),
    .io_data_out_b_field_type_26_sub_class_id(meta_table_io_data_out_b_field_type_26_sub_class_id),
    .io_data_out_b_field_type_27_is_repeated(meta_table_io_data_out_b_field_type_27_is_repeated),
    .io_data_out_b_field_type_27_field_type(meta_table_io_data_out_b_field_type_27_field_type),
    .io_data_out_b_field_type_27_sub_class_id(meta_table_io_data_out_b_field_type_27_sub_class_id),
    .io_data_out_b_field_type_28_is_repeated(meta_table_io_data_out_b_field_type_28_is_repeated),
    .io_data_out_b_field_type_28_field_type(meta_table_io_data_out_b_field_type_28_field_type),
    .io_data_out_b_field_type_28_sub_class_id(meta_table_io_data_out_b_field_type_28_sub_class_id),
    .io_data_out_b_field_type_29_is_repeated(meta_table_io_data_out_b_field_type_29_is_repeated),
    .io_data_out_b_field_type_29_field_type(meta_table_io_data_out_b_field_type_29_field_type),
    .io_data_out_b_field_type_29_sub_class_id(meta_table_io_data_out_b_field_type_29_sub_class_id),
    .io_data_out_b_field_type_30_is_repeated(meta_table_io_data_out_b_field_type_30_is_repeated),
    .io_data_out_b_field_type_30_field_type(meta_table_io_data_out_b_field_type_30_field_type),
    .io_data_out_b_field_type_30_sub_class_id(meta_table_io_data_out_b_field_type_30_sub_class_id),
    .io_data_out_b_field_type_31_is_repeated(meta_table_io_data_out_b_field_type_31_is_repeated),
    .io_data_out_b_field_type_31_field_type(meta_table_io_data_out_b_field_type_31_field_type),
    .io_data_out_b_field_type_31_sub_class_id(meta_table_io_data_out_b_field_type_31_sub_class_id),
    .io_data_out_b_field_type_32_is_repeated(meta_table_io_data_out_b_field_type_32_is_repeated),
    .io_data_out_b_field_type_32_field_type(meta_table_io_data_out_b_field_type_32_field_type),
    .io_data_out_b_field_type_32_sub_class_id(meta_table_io_data_out_b_field_type_32_sub_class_id)
  );
  assign io_class_meta_init_ready = 1'h1; // @[ClassMetaTable.scala 76:48]
  assign io_s_class_meta_req_ready = s_class_meta_req_fifo_io_in_ready; // @[ClassMetaTable.scala 56:47]
  assign io_s_class_meta_rsp_valid = state == 2'h1; // @[ClassMetaTable.scala 104:16]
  assign io_s_class_meta_rsp_bits_class_meta_max_field_num = state == 2'h1 ? meta_table_io_data_out_b_max_field_num : 8'h0
    ; // @[ClassMetaTable.scala 104:26 ClassMetaTable.scala 107:51 Util.scala 13:25]
  assign io_s_class_meta_rsp_bits_class_meta_field_type_0_is_repeated = state == 2'h1 &
    meta_table_io_data_out_b_field_type_0_is_repeated; // @[ClassMetaTable.scala 104:26 ClassMetaTable.scala 107:51 Util.scala 13:25]
  assign io_s_class_meta_rsp_bits_class_meta_field_type_0_field_type = state == 2'h1 ?
    meta_table_io_data_out_b_field_type_0_field_type : 5'h0; // @[ClassMetaTable.scala 104:26 ClassMetaTable.scala 107:51 Util.scala 13:25]
  assign io_s_class_meta_rsp_bits_class_meta_field_type_0_sub_class_id = state == 2'h1 ?
    meta_table_io_data_out_b_field_type_0_sub_class_id : 16'h0; // @[ClassMetaTable.scala 104:26 ClassMetaTable.scala 107:51 Util.scala 13:25]
  assign io_s_class_meta_rsp_bits_class_meta_field_type_1_is_repeated = state == 2'h1 &
    meta_table_io_data_out_b_field_type_1_is_repeated; // @[ClassMetaTable.scala 104:26 ClassMetaTable.scala 107:51 Util.scala 13:25]
  assign io_s_class_meta_rsp_bits_class_meta_field_type_1_field_type = state == 2'h1 ?
    meta_table_io_data_out_b_field_type_1_field_type : 5'h0; // @[ClassMetaTable.scala 104:26 ClassMetaTable.scala 107:51 Util.scala 13:25]
  assign io_s_class_meta_rsp_bits_class_meta_field_type_1_sub_class_id = state == 2'h1 ?
    meta_table_io_data_out_b_field_type_1_sub_class_id : 16'h0; // @[ClassMetaTable.scala 104:26 ClassMetaTable.scala 107:51 Util.scala 13:25]
  assign io_s_class_meta_rsp_bits_class_meta_field_type_2_is_repeated = state == 2'h1 &
    meta_table_io_data_out_b_field_type_2_is_repeated; // @[ClassMetaTable.scala 104:26 ClassMetaTable.scala 107:51 Util.scala 13:25]
  assign io_s_class_meta_rsp_bits_class_meta_field_type_2_field_type = state == 2'h1 ?
    meta_table_io_data_out_b_field_type_2_field_type : 5'h0; // @[ClassMetaTable.scala 104:26 ClassMetaTable.scala 107:51 Util.scala 13:25]
  assign io_s_class_meta_rsp_bits_class_meta_field_type_2_sub_class_id = state == 2'h1 ?
    meta_table_io_data_out_b_field_type_2_sub_class_id : 16'h0; // @[ClassMetaTable.scala 104:26 ClassMetaTable.scala 107:51 Util.scala 13:25]
  assign io_s_class_meta_rsp_bits_class_meta_field_type_3_is_repeated = state == 2'h1 &
    meta_table_io_data_out_b_field_type_3_is_repeated; // @[ClassMetaTable.scala 104:26 ClassMetaTable.scala 107:51 Util.scala 13:25]
  assign io_s_class_meta_rsp_bits_class_meta_field_type_3_field_type = state == 2'h1 ?
    meta_table_io_data_out_b_field_type_3_field_type : 5'h0; // @[ClassMetaTable.scala 104:26 ClassMetaTable.scala 107:51 Util.scala 13:25]
  assign io_s_class_meta_rsp_bits_class_meta_field_type_3_sub_class_id = state == 2'h1 ?
    meta_table_io_data_out_b_field_type_3_sub_class_id : 16'h0; // @[ClassMetaTable.scala 104:26 ClassMetaTable.scala 107:51 Util.scala 13:25]
  assign io_s_class_meta_rsp_bits_class_meta_field_type_4_is_repeated = state == 2'h1 &
    meta_table_io_data_out_b_field_type_4_is_repeated; // @[ClassMetaTable.scala 104:26 ClassMetaTable.scala 107:51 Util.scala 13:25]
  assign io_s_class_meta_rsp_bits_class_meta_field_type_4_field_type = state == 2'h1 ?
    meta_table_io_data_out_b_field_type_4_field_type : 5'h0; // @[ClassMetaTable.scala 104:26 ClassMetaTable.scala 107:51 Util.scala 13:25]
  assign io_s_class_meta_rsp_bits_class_meta_field_type_4_sub_class_id = state == 2'h1 ?
    meta_table_io_data_out_b_field_type_4_sub_class_id : 16'h0; // @[ClassMetaTable.scala 104:26 ClassMetaTable.scala 107:51 Util.scala 13:25]
  assign io_s_class_meta_rsp_bits_class_meta_field_type_5_is_repeated = state == 2'h1 &
    meta_table_io_data_out_b_field_type_5_is_repeated; // @[ClassMetaTable.scala 104:26 ClassMetaTable.scala 107:51 Util.scala 13:25]
  assign io_s_class_meta_rsp_bits_class_meta_field_type_5_field_type = state == 2'h1 ?
    meta_table_io_data_out_b_field_type_5_field_type : 5'h0; // @[ClassMetaTable.scala 104:26 ClassMetaTable.scala 107:51 Util.scala 13:25]
  assign io_s_class_meta_rsp_bits_class_meta_field_type_5_sub_class_id = state == 2'h1 ?
    meta_table_io_data_out_b_field_type_5_sub_class_id : 16'h0; // @[ClassMetaTable.scala 104:26 ClassMetaTable.scala 107:51 Util.scala 13:25]
  assign io_s_class_meta_rsp_bits_class_meta_field_type_6_is_repeated = state == 2'h1 &
    meta_table_io_data_out_b_field_type_6_is_repeated; // @[ClassMetaTable.scala 104:26 ClassMetaTable.scala 107:51 Util.scala 13:25]
  assign io_s_class_meta_rsp_bits_class_meta_field_type_6_field_type = state == 2'h1 ?
    meta_table_io_data_out_b_field_type_6_field_type : 5'h0; // @[ClassMetaTable.scala 104:26 ClassMetaTable.scala 107:51 Util.scala 13:25]
  assign io_s_class_meta_rsp_bits_class_meta_field_type_6_sub_class_id = state == 2'h1 ?
    meta_table_io_data_out_b_field_type_6_sub_class_id : 16'h0; // @[ClassMetaTable.scala 104:26 ClassMetaTable.scala 107:51 Util.scala 13:25]
  assign io_s_class_meta_rsp_bits_class_meta_field_type_7_is_repeated = state == 2'h1 &
    meta_table_io_data_out_b_field_type_7_is_repeated; // @[ClassMetaTable.scala 104:26 ClassMetaTable.scala 107:51 Util.scala 13:25]
  assign io_s_class_meta_rsp_bits_class_meta_field_type_7_field_type = state == 2'h1 ?
    meta_table_io_data_out_b_field_type_7_field_type : 5'h0; // @[ClassMetaTable.scala 104:26 ClassMetaTable.scala 107:51 Util.scala 13:25]
  assign io_s_class_meta_rsp_bits_class_meta_field_type_7_sub_class_id = state == 2'h1 ?
    meta_table_io_data_out_b_field_type_7_sub_class_id : 16'h0; // @[ClassMetaTable.scala 104:26 ClassMetaTable.scala 107:51 Util.scala 13:25]
  assign io_s_class_meta_rsp_bits_class_meta_field_type_8_is_repeated = state == 2'h1 &
    meta_table_io_data_out_b_field_type_8_is_repeated; // @[ClassMetaTable.scala 104:26 ClassMetaTable.scala 107:51 Util.scala 13:25]
  assign io_s_class_meta_rsp_bits_class_meta_field_type_8_field_type = state == 2'h1 ?
    meta_table_io_data_out_b_field_type_8_field_type : 5'h0; // @[ClassMetaTable.scala 104:26 ClassMetaTable.scala 107:51 Util.scala 13:25]
  assign io_s_class_meta_rsp_bits_class_meta_field_type_8_sub_class_id = state == 2'h1 ?
    meta_table_io_data_out_b_field_type_8_sub_class_id : 16'h0; // @[ClassMetaTable.scala 104:26 ClassMetaTable.scala 107:51 Util.scala 13:25]
  assign io_s_class_meta_rsp_bits_class_meta_field_type_9_is_repeated = state == 2'h1 &
    meta_table_io_data_out_b_field_type_9_is_repeated; // @[ClassMetaTable.scala 104:26 ClassMetaTable.scala 107:51 Util.scala 13:25]
  assign io_s_class_meta_rsp_bits_class_meta_field_type_9_field_type = state == 2'h1 ?
    meta_table_io_data_out_b_field_type_9_field_type : 5'h0; // @[ClassMetaTable.scala 104:26 ClassMetaTable.scala 107:51 Util.scala 13:25]
  assign io_s_class_meta_rsp_bits_class_meta_field_type_9_sub_class_id = state == 2'h1 ?
    meta_table_io_data_out_b_field_type_9_sub_class_id : 16'h0; // @[ClassMetaTable.scala 104:26 ClassMetaTable.scala 107:51 Util.scala 13:25]
  assign io_s_class_meta_rsp_bits_class_meta_field_type_10_is_repeated = state == 2'h1 &
    meta_table_io_data_out_b_field_type_10_is_repeated; // @[ClassMetaTable.scala 104:26 ClassMetaTable.scala 107:51 Util.scala 13:25]
  assign io_s_class_meta_rsp_bits_class_meta_field_type_10_field_type = state == 2'h1 ?
    meta_table_io_data_out_b_field_type_10_field_type : 5'h0; // @[ClassMetaTable.scala 104:26 ClassMetaTable.scala 107:51 Util.scala 13:25]
  assign io_s_class_meta_rsp_bits_class_meta_field_type_10_sub_class_id = state == 2'h1 ?
    meta_table_io_data_out_b_field_type_10_sub_class_id : 16'h0; // @[ClassMetaTable.scala 104:26 ClassMetaTable.scala 107:51 Util.scala 13:25]
  assign io_s_class_meta_rsp_bits_class_meta_field_type_11_is_repeated = state == 2'h1 &
    meta_table_io_data_out_b_field_type_11_is_repeated; // @[ClassMetaTable.scala 104:26 ClassMetaTable.scala 107:51 Util.scala 13:25]
  assign io_s_class_meta_rsp_bits_class_meta_field_type_11_field_type = state == 2'h1 ?
    meta_table_io_data_out_b_field_type_11_field_type : 5'h0; // @[ClassMetaTable.scala 104:26 ClassMetaTable.scala 107:51 Util.scala 13:25]
  assign io_s_class_meta_rsp_bits_class_meta_field_type_11_sub_class_id = state == 2'h1 ?
    meta_table_io_data_out_b_field_type_11_sub_class_id : 16'h0; // @[ClassMetaTable.scala 104:26 ClassMetaTable.scala 107:51 Util.scala 13:25]
  assign io_s_class_meta_rsp_bits_class_meta_field_type_12_is_repeated = state == 2'h1 &
    meta_table_io_data_out_b_field_type_12_is_repeated; // @[ClassMetaTable.scala 104:26 ClassMetaTable.scala 107:51 Util.scala 13:25]
  assign io_s_class_meta_rsp_bits_class_meta_field_type_12_field_type = state == 2'h1 ?
    meta_table_io_data_out_b_field_type_12_field_type : 5'h0; // @[ClassMetaTable.scala 104:26 ClassMetaTable.scala 107:51 Util.scala 13:25]
  assign io_s_class_meta_rsp_bits_class_meta_field_type_12_sub_class_id = state == 2'h1 ?
    meta_table_io_data_out_b_field_type_12_sub_class_id : 16'h0; // @[ClassMetaTable.scala 104:26 ClassMetaTable.scala 107:51 Util.scala 13:25]
  assign io_s_class_meta_rsp_bits_class_meta_field_type_13_is_repeated = state == 2'h1 &
    meta_table_io_data_out_b_field_type_13_is_repeated; // @[ClassMetaTable.scala 104:26 ClassMetaTable.scala 107:51 Util.scala 13:25]
  assign io_s_class_meta_rsp_bits_class_meta_field_type_13_field_type = state == 2'h1 ?
    meta_table_io_data_out_b_field_type_13_field_type : 5'h0; // @[ClassMetaTable.scala 104:26 ClassMetaTable.scala 107:51 Util.scala 13:25]
  assign io_s_class_meta_rsp_bits_class_meta_field_type_13_sub_class_id = state == 2'h1 ?
    meta_table_io_data_out_b_field_type_13_sub_class_id : 16'h0; // @[ClassMetaTable.scala 104:26 ClassMetaTable.scala 107:51 Util.scala 13:25]
  assign io_s_class_meta_rsp_bits_class_meta_field_type_14_is_repeated = state == 2'h1 &
    meta_table_io_data_out_b_field_type_14_is_repeated; // @[ClassMetaTable.scala 104:26 ClassMetaTable.scala 107:51 Util.scala 13:25]
  assign io_s_class_meta_rsp_bits_class_meta_field_type_14_field_type = state == 2'h1 ?
    meta_table_io_data_out_b_field_type_14_field_type : 5'h0; // @[ClassMetaTable.scala 104:26 ClassMetaTable.scala 107:51 Util.scala 13:25]
  assign io_s_class_meta_rsp_bits_class_meta_field_type_14_sub_class_id = state == 2'h1 ?
    meta_table_io_data_out_b_field_type_14_sub_class_id : 16'h0; // @[ClassMetaTable.scala 104:26 ClassMetaTable.scala 107:51 Util.scala 13:25]
  assign io_s_class_meta_rsp_bits_class_meta_field_type_15_is_repeated = state == 2'h1 &
    meta_table_io_data_out_b_field_type_15_is_repeated; // @[ClassMetaTable.scala 104:26 ClassMetaTable.scala 107:51 Util.scala 13:25]
  assign io_s_class_meta_rsp_bits_class_meta_field_type_15_field_type = state == 2'h1 ?
    meta_table_io_data_out_b_field_type_15_field_type : 5'h0; // @[ClassMetaTable.scala 104:26 ClassMetaTable.scala 107:51 Util.scala 13:25]
  assign io_s_class_meta_rsp_bits_class_meta_field_type_15_sub_class_id = state == 2'h1 ?
    meta_table_io_data_out_b_field_type_15_sub_class_id : 16'h0; // @[ClassMetaTable.scala 104:26 ClassMetaTable.scala 107:51 Util.scala 13:25]
  assign io_s_class_meta_rsp_bits_class_meta_field_type_16_is_repeated = state == 2'h1 &
    meta_table_io_data_out_b_field_type_16_is_repeated; // @[ClassMetaTable.scala 104:26 ClassMetaTable.scala 107:51 Util.scala 13:25]
  assign io_s_class_meta_rsp_bits_class_meta_field_type_16_field_type = state == 2'h1 ?
    meta_table_io_data_out_b_field_type_16_field_type : 5'h0; // @[ClassMetaTable.scala 104:26 ClassMetaTable.scala 107:51 Util.scala 13:25]
  assign io_s_class_meta_rsp_bits_class_meta_field_type_16_sub_class_id = state == 2'h1 ?
    meta_table_io_data_out_b_field_type_16_sub_class_id : 16'h0; // @[ClassMetaTable.scala 104:26 ClassMetaTable.scala 107:51 Util.scala 13:25]
  assign io_s_class_meta_rsp_bits_class_meta_field_type_17_is_repeated = state == 2'h1 &
    meta_table_io_data_out_b_field_type_17_is_repeated; // @[ClassMetaTable.scala 104:26 ClassMetaTable.scala 107:51 Util.scala 13:25]
  assign io_s_class_meta_rsp_bits_class_meta_field_type_17_field_type = state == 2'h1 ?
    meta_table_io_data_out_b_field_type_17_field_type : 5'h0; // @[ClassMetaTable.scala 104:26 ClassMetaTable.scala 107:51 Util.scala 13:25]
  assign io_s_class_meta_rsp_bits_class_meta_field_type_17_sub_class_id = state == 2'h1 ?
    meta_table_io_data_out_b_field_type_17_sub_class_id : 16'h0; // @[ClassMetaTable.scala 104:26 ClassMetaTable.scala 107:51 Util.scala 13:25]
  assign io_s_class_meta_rsp_bits_class_meta_field_type_18_is_repeated = state == 2'h1 &
    meta_table_io_data_out_b_field_type_18_is_repeated; // @[ClassMetaTable.scala 104:26 ClassMetaTable.scala 107:51 Util.scala 13:25]
  assign io_s_class_meta_rsp_bits_class_meta_field_type_18_field_type = state == 2'h1 ?
    meta_table_io_data_out_b_field_type_18_field_type : 5'h0; // @[ClassMetaTable.scala 104:26 ClassMetaTable.scala 107:51 Util.scala 13:25]
  assign io_s_class_meta_rsp_bits_class_meta_field_type_18_sub_class_id = state == 2'h1 ?
    meta_table_io_data_out_b_field_type_18_sub_class_id : 16'h0; // @[ClassMetaTable.scala 104:26 ClassMetaTable.scala 107:51 Util.scala 13:25]
  assign io_s_class_meta_rsp_bits_class_meta_field_type_19_is_repeated = state == 2'h1 &
    meta_table_io_data_out_b_field_type_19_is_repeated; // @[ClassMetaTable.scala 104:26 ClassMetaTable.scala 107:51 Util.scala 13:25]
  assign io_s_class_meta_rsp_bits_class_meta_field_type_19_field_type = state == 2'h1 ?
    meta_table_io_data_out_b_field_type_19_field_type : 5'h0; // @[ClassMetaTable.scala 104:26 ClassMetaTable.scala 107:51 Util.scala 13:25]
  assign io_s_class_meta_rsp_bits_class_meta_field_type_19_sub_class_id = state == 2'h1 ?
    meta_table_io_data_out_b_field_type_19_sub_class_id : 16'h0; // @[ClassMetaTable.scala 104:26 ClassMetaTable.scala 107:51 Util.scala 13:25]
  assign io_s_class_meta_rsp_bits_class_meta_field_type_20_is_repeated = state == 2'h1 &
    meta_table_io_data_out_b_field_type_20_is_repeated; // @[ClassMetaTable.scala 104:26 ClassMetaTable.scala 107:51 Util.scala 13:25]
  assign io_s_class_meta_rsp_bits_class_meta_field_type_20_field_type = state == 2'h1 ?
    meta_table_io_data_out_b_field_type_20_field_type : 5'h0; // @[ClassMetaTable.scala 104:26 ClassMetaTable.scala 107:51 Util.scala 13:25]
  assign io_s_class_meta_rsp_bits_class_meta_field_type_20_sub_class_id = state == 2'h1 ?
    meta_table_io_data_out_b_field_type_20_sub_class_id : 16'h0; // @[ClassMetaTable.scala 104:26 ClassMetaTable.scala 107:51 Util.scala 13:25]
  assign io_s_class_meta_rsp_bits_class_meta_field_type_21_is_repeated = state == 2'h1 &
    meta_table_io_data_out_b_field_type_21_is_repeated; // @[ClassMetaTable.scala 104:26 ClassMetaTable.scala 107:51 Util.scala 13:25]
  assign io_s_class_meta_rsp_bits_class_meta_field_type_21_field_type = state == 2'h1 ?
    meta_table_io_data_out_b_field_type_21_field_type : 5'h0; // @[ClassMetaTable.scala 104:26 ClassMetaTable.scala 107:51 Util.scala 13:25]
  assign io_s_class_meta_rsp_bits_class_meta_field_type_21_sub_class_id = state == 2'h1 ?
    meta_table_io_data_out_b_field_type_21_sub_class_id : 16'h0; // @[ClassMetaTable.scala 104:26 ClassMetaTable.scala 107:51 Util.scala 13:25]
  assign io_s_class_meta_rsp_bits_class_meta_field_type_22_is_repeated = state == 2'h1 &
    meta_table_io_data_out_b_field_type_22_is_repeated; // @[ClassMetaTable.scala 104:26 ClassMetaTable.scala 107:51 Util.scala 13:25]
  assign io_s_class_meta_rsp_bits_class_meta_field_type_22_field_type = state == 2'h1 ?
    meta_table_io_data_out_b_field_type_22_field_type : 5'h0; // @[ClassMetaTable.scala 104:26 ClassMetaTable.scala 107:51 Util.scala 13:25]
  assign io_s_class_meta_rsp_bits_class_meta_field_type_22_sub_class_id = state == 2'h1 ?
    meta_table_io_data_out_b_field_type_22_sub_class_id : 16'h0; // @[ClassMetaTable.scala 104:26 ClassMetaTable.scala 107:51 Util.scala 13:25]
  assign io_s_class_meta_rsp_bits_class_meta_field_type_23_is_repeated = state == 2'h1 &
    meta_table_io_data_out_b_field_type_23_is_repeated; // @[ClassMetaTable.scala 104:26 ClassMetaTable.scala 107:51 Util.scala 13:25]
  assign io_s_class_meta_rsp_bits_class_meta_field_type_23_field_type = state == 2'h1 ?
    meta_table_io_data_out_b_field_type_23_field_type : 5'h0; // @[ClassMetaTable.scala 104:26 ClassMetaTable.scala 107:51 Util.scala 13:25]
  assign io_s_class_meta_rsp_bits_class_meta_field_type_23_sub_class_id = state == 2'h1 ?
    meta_table_io_data_out_b_field_type_23_sub_class_id : 16'h0; // @[ClassMetaTable.scala 104:26 ClassMetaTable.scala 107:51 Util.scala 13:25]
  assign io_s_class_meta_rsp_bits_class_meta_field_type_24_is_repeated = state == 2'h1 &
    meta_table_io_data_out_b_field_type_24_is_repeated; // @[ClassMetaTable.scala 104:26 ClassMetaTable.scala 107:51 Util.scala 13:25]
  assign io_s_class_meta_rsp_bits_class_meta_field_type_24_field_type = state == 2'h1 ?
    meta_table_io_data_out_b_field_type_24_field_type : 5'h0; // @[ClassMetaTable.scala 104:26 ClassMetaTable.scala 107:51 Util.scala 13:25]
  assign io_s_class_meta_rsp_bits_class_meta_field_type_24_sub_class_id = state == 2'h1 ?
    meta_table_io_data_out_b_field_type_24_sub_class_id : 16'h0; // @[ClassMetaTable.scala 104:26 ClassMetaTable.scala 107:51 Util.scala 13:25]
  assign io_s_class_meta_rsp_bits_class_meta_field_type_25_is_repeated = state == 2'h1 &
    meta_table_io_data_out_b_field_type_25_is_repeated; // @[ClassMetaTable.scala 104:26 ClassMetaTable.scala 107:51 Util.scala 13:25]
  assign io_s_class_meta_rsp_bits_class_meta_field_type_25_field_type = state == 2'h1 ?
    meta_table_io_data_out_b_field_type_25_field_type : 5'h0; // @[ClassMetaTable.scala 104:26 ClassMetaTable.scala 107:51 Util.scala 13:25]
  assign io_s_class_meta_rsp_bits_class_meta_field_type_25_sub_class_id = state == 2'h1 ?
    meta_table_io_data_out_b_field_type_25_sub_class_id : 16'h0; // @[ClassMetaTable.scala 104:26 ClassMetaTable.scala 107:51 Util.scala 13:25]
  assign io_s_class_meta_rsp_bits_class_meta_field_type_26_is_repeated = state == 2'h1 &
    meta_table_io_data_out_b_field_type_26_is_repeated; // @[ClassMetaTable.scala 104:26 ClassMetaTable.scala 107:51 Util.scala 13:25]
  assign io_s_class_meta_rsp_bits_class_meta_field_type_26_field_type = state == 2'h1 ?
    meta_table_io_data_out_b_field_type_26_field_type : 5'h0; // @[ClassMetaTable.scala 104:26 ClassMetaTable.scala 107:51 Util.scala 13:25]
  assign io_s_class_meta_rsp_bits_class_meta_field_type_26_sub_class_id = state == 2'h1 ?
    meta_table_io_data_out_b_field_type_26_sub_class_id : 16'h0; // @[ClassMetaTable.scala 104:26 ClassMetaTable.scala 107:51 Util.scala 13:25]
  assign io_s_class_meta_rsp_bits_class_meta_field_type_27_is_repeated = state == 2'h1 &
    meta_table_io_data_out_b_field_type_27_is_repeated; // @[ClassMetaTable.scala 104:26 ClassMetaTable.scala 107:51 Util.scala 13:25]
  assign io_s_class_meta_rsp_bits_class_meta_field_type_27_field_type = state == 2'h1 ?
    meta_table_io_data_out_b_field_type_27_field_type : 5'h0; // @[ClassMetaTable.scala 104:26 ClassMetaTable.scala 107:51 Util.scala 13:25]
  assign io_s_class_meta_rsp_bits_class_meta_field_type_27_sub_class_id = state == 2'h1 ?
    meta_table_io_data_out_b_field_type_27_sub_class_id : 16'h0; // @[ClassMetaTable.scala 104:26 ClassMetaTable.scala 107:51 Util.scala 13:25]
  assign io_s_class_meta_rsp_bits_class_meta_field_type_28_is_repeated = state == 2'h1 &
    meta_table_io_data_out_b_field_type_28_is_repeated; // @[ClassMetaTable.scala 104:26 ClassMetaTable.scala 107:51 Util.scala 13:25]
  assign io_s_class_meta_rsp_bits_class_meta_field_type_28_field_type = state == 2'h1 ?
    meta_table_io_data_out_b_field_type_28_field_type : 5'h0; // @[ClassMetaTable.scala 104:26 ClassMetaTable.scala 107:51 Util.scala 13:25]
  assign io_s_class_meta_rsp_bits_class_meta_field_type_28_sub_class_id = state == 2'h1 ?
    meta_table_io_data_out_b_field_type_28_sub_class_id : 16'h0; // @[ClassMetaTable.scala 104:26 ClassMetaTable.scala 107:51 Util.scala 13:25]
  assign io_s_class_meta_rsp_bits_class_meta_field_type_29_is_repeated = state == 2'h1 &
    meta_table_io_data_out_b_field_type_29_is_repeated; // @[ClassMetaTable.scala 104:26 ClassMetaTable.scala 107:51 Util.scala 13:25]
  assign io_s_class_meta_rsp_bits_class_meta_field_type_29_field_type = state == 2'h1 ?
    meta_table_io_data_out_b_field_type_29_field_type : 5'h0; // @[ClassMetaTable.scala 104:26 ClassMetaTable.scala 107:51 Util.scala 13:25]
  assign io_s_class_meta_rsp_bits_class_meta_field_type_29_sub_class_id = state == 2'h1 ?
    meta_table_io_data_out_b_field_type_29_sub_class_id : 16'h0; // @[ClassMetaTable.scala 104:26 ClassMetaTable.scala 107:51 Util.scala 13:25]
  assign io_s_class_meta_rsp_bits_class_meta_field_type_30_is_repeated = state == 2'h1 &
    meta_table_io_data_out_b_field_type_30_is_repeated; // @[ClassMetaTable.scala 104:26 ClassMetaTable.scala 107:51 Util.scala 13:25]
  assign io_s_class_meta_rsp_bits_class_meta_field_type_30_field_type = state == 2'h1 ?
    meta_table_io_data_out_b_field_type_30_field_type : 5'h0; // @[ClassMetaTable.scala 104:26 ClassMetaTable.scala 107:51 Util.scala 13:25]
  assign io_s_class_meta_rsp_bits_class_meta_field_type_30_sub_class_id = state == 2'h1 ?
    meta_table_io_data_out_b_field_type_30_sub_class_id : 16'h0; // @[ClassMetaTable.scala 104:26 ClassMetaTable.scala 107:51 Util.scala 13:25]
  assign io_s_class_meta_rsp_bits_class_meta_field_type_31_is_repeated = state == 2'h1 &
    meta_table_io_data_out_b_field_type_31_is_repeated; // @[ClassMetaTable.scala 104:26 ClassMetaTable.scala 107:51 Util.scala 13:25]
  assign io_s_class_meta_rsp_bits_class_meta_field_type_31_field_type = state == 2'h1 ?
    meta_table_io_data_out_b_field_type_31_field_type : 5'h0; // @[ClassMetaTable.scala 104:26 ClassMetaTable.scala 107:51 Util.scala 13:25]
  assign io_s_class_meta_rsp_bits_class_meta_field_type_31_sub_class_id = state == 2'h1 ?
    meta_table_io_data_out_b_field_type_31_sub_class_id : 16'h0; // @[ClassMetaTable.scala 104:26 ClassMetaTable.scala 107:51 Util.scala 13:25]
  assign io_s_class_meta_rsp_bits_class_meta_field_type_32_is_repeated = state == 2'h1 &
    meta_table_io_data_out_b_field_type_32_is_repeated; // @[ClassMetaTable.scala 104:26 ClassMetaTable.scala 107:51 Util.scala 13:25]
  assign io_s_class_meta_rsp_bits_class_meta_field_type_32_field_type = state == 2'h1 ?
    meta_table_io_data_out_b_field_type_32_field_type : 5'h0; // @[ClassMetaTable.scala 104:26 ClassMetaTable.scala 107:51 Util.scala 13:25]
  assign io_s_class_meta_rsp_bits_class_meta_field_type_32_sub_class_id = state == 2'h1 ?
    meta_table_io_data_out_b_field_type_32_sub_class_id : 16'h0; // @[ClassMetaTable.scala 104:26 ClassMetaTable.scala 107:51 Util.scala 13:25]
  assign counter_5 = counter;
  assign s_class_meta_req_fifo_clock = clock;
  assign s_class_meta_req_fifo_reset = reset;
  assign s_class_meta_req_fifo_io_in_valid = io_s_class_meta_req_valid; // @[ClassMetaTable.scala 56:47]
  assign s_class_meta_req_fifo_io_in_bits_class_id = io_s_class_meta_req_bits_class_id; // @[ClassMetaTable.scala 56:47]
  assign s_class_meta_req_fifo_io_out_ready = ~io_class_meta_init_valid & state == 2'h0; // @[ClassMetaTable.scala 74:88]
  assign d_class_meta_req_fifo_clock = clock;
  assign d_class_meta_req_fifo_reset = reset;
  assign d_class_meta_req_fifo_io_in_valid = 1'h0; // @[ClassMetaTable.scala 57:47]
  assign d_class_meta_req_fifo_io_in_bits_class_id = 10'h0; // @[ClassMetaTable.scala 57:47]
  assign d_class_meta_req_fifo_io_out_ready = _s_class_meta_req_fifo_io_out_ready_T_1 & ~
    s_class_meta_req_fifo_io_out_valid & _s_class_meta_req_fifo_io_out_ready_T_2; // @[ClassMetaTable.scala 75:135]
  assign meta_table_clock = clock;
  assign meta_table_reset = reset;
  assign meta_table_io_addr_a = _T ? io_class_meta_init_bits_class_id : 10'h0; // @[ClassMetaTable.scala 85:36 ClassMetaTable.scala 86:49 ClassMetaTable.scala 69:42]
  assign meta_table_io_addr_b = _T ? 10'h0 : _GEN_4; // @[ClassMetaTable.scala 85:36 ClassMetaTable.scala 70:42]
  assign meta_table_io_wr_en_a = io_class_meta_init_ready & io_class_meta_init_valid; // @[Decoupled.scala 40:37]
  assign meta_table_io_data_in_a_class_length = _T ? io_class_meta_init_bits_desc_state_class_length : 16'h0; // @[ClassMetaTable.scala 85:36 ClassMetaTable.scala 88:49 ClassMetaTable.scala 72:42]
  assign meta_table_io_data_in_a_max_field_num = _T ? io_class_meta_init_bits_desc_state_max_field_num : 8'h0; // @[ClassMetaTable.scala 85:36 ClassMetaTable.scala 88:49 ClassMetaTable.scala 72:42]
  assign meta_table_io_data_in_a_field_type_0_is_repeated = _T &
    io_class_meta_init_bits_desc_state_field_type_0_is_repeated; // @[ClassMetaTable.scala 85:36 ClassMetaTable.scala 88:49 ClassMetaTable.scala 72:42]
  assign meta_table_io_data_in_a_field_type_0_field_type = _T ?
    io_class_meta_init_bits_desc_state_field_type_0_field_type : 5'h0; // @[ClassMetaTable.scala 85:36 ClassMetaTable.scala 88:49 ClassMetaTable.scala 72:42]
  assign meta_table_io_data_in_a_field_type_0_sub_class_id = _T ?
    io_class_meta_init_bits_desc_state_field_type_0_sub_class_id : 16'h0; // @[ClassMetaTable.scala 85:36 ClassMetaTable.scala 88:49 ClassMetaTable.scala 72:42]
  assign meta_table_io_data_in_a_field_type_0_is_host = _T & io_class_meta_init_bits_desc_state_field_type_0_is_host; // @[ClassMetaTable.scala 85:36 ClassMetaTable.scala 88:49 ClassMetaTable.scala 72:42]
  assign meta_table_io_data_in_a_field_type_1_is_repeated = _T &
    io_class_meta_init_bits_desc_state_field_type_1_is_repeated; // @[ClassMetaTable.scala 85:36 ClassMetaTable.scala 88:49 ClassMetaTable.scala 72:42]
  assign meta_table_io_data_in_a_field_type_1_field_type = _T ?
    io_class_meta_init_bits_desc_state_field_type_1_field_type : 5'h0; // @[ClassMetaTable.scala 85:36 ClassMetaTable.scala 88:49 ClassMetaTable.scala 72:42]
  assign meta_table_io_data_in_a_field_type_1_sub_class_id = _T ?
    io_class_meta_init_bits_desc_state_field_type_1_sub_class_id : 16'h0; // @[ClassMetaTable.scala 85:36 ClassMetaTable.scala 88:49 ClassMetaTable.scala 72:42]
  assign meta_table_io_data_in_a_field_type_1_is_host = _T & io_class_meta_init_bits_desc_state_field_type_1_is_host; // @[ClassMetaTable.scala 85:36 ClassMetaTable.scala 88:49 ClassMetaTable.scala 72:42]
  assign meta_table_io_data_in_a_field_type_2_is_repeated = _T &
    io_class_meta_init_bits_desc_state_field_type_2_is_repeated; // @[ClassMetaTable.scala 85:36 ClassMetaTable.scala 88:49 ClassMetaTable.scala 72:42]
  assign meta_table_io_data_in_a_field_type_2_field_type = _T ?
    io_class_meta_init_bits_desc_state_field_type_2_field_type : 5'h0; // @[ClassMetaTable.scala 85:36 ClassMetaTable.scala 88:49 ClassMetaTable.scala 72:42]
  assign meta_table_io_data_in_a_field_type_2_sub_class_id = _T ?
    io_class_meta_init_bits_desc_state_field_type_2_sub_class_id : 16'h0; // @[ClassMetaTable.scala 85:36 ClassMetaTable.scala 88:49 ClassMetaTable.scala 72:42]
  assign meta_table_io_data_in_a_field_type_2_is_host = _T & io_class_meta_init_bits_desc_state_field_type_2_is_host; // @[ClassMetaTable.scala 85:36 ClassMetaTable.scala 88:49 ClassMetaTable.scala 72:42]
  assign meta_table_io_data_in_a_field_type_3_is_repeated = _T &
    io_class_meta_init_bits_desc_state_field_type_3_is_repeated; // @[ClassMetaTable.scala 85:36 ClassMetaTable.scala 88:49 ClassMetaTable.scala 72:42]
  assign meta_table_io_data_in_a_field_type_3_field_type = _T ?
    io_class_meta_init_bits_desc_state_field_type_3_field_type : 5'h0; // @[ClassMetaTable.scala 85:36 ClassMetaTable.scala 88:49 ClassMetaTable.scala 72:42]
  assign meta_table_io_data_in_a_field_type_3_sub_class_id = _T ?
    io_class_meta_init_bits_desc_state_field_type_3_sub_class_id : 16'h0; // @[ClassMetaTable.scala 85:36 ClassMetaTable.scala 88:49 ClassMetaTable.scala 72:42]
  assign meta_table_io_data_in_a_field_type_3_is_host = _T & io_class_meta_init_bits_desc_state_field_type_3_is_host; // @[ClassMetaTable.scala 85:36 ClassMetaTable.scala 88:49 ClassMetaTable.scala 72:42]
  assign meta_table_io_data_in_a_field_type_4_is_repeated = _T &
    io_class_meta_init_bits_desc_state_field_type_4_is_repeated; // @[ClassMetaTable.scala 85:36 ClassMetaTable.scala 88:49 ClassMetaTable.scala 72:42]
  assign meta_table_io_data_in_a_field_type_4_field_type = _T ?
    io_class_meta_init_bits_desc_state_field_type_4_field_type : 5'h0; // @[ClassMetaTable.scala 85:36 ClassMetaTable.scala 88:49 ClassMetaTable.scala 72:42]
  assign meta_table_io_data_in_a_field_type_4_sub_class_id = _T ?
    io_class_meta_init_bits_desc_state_field_type_4_sub_class_id : 16'h0; // @[ClassMetaTable.scala 85:36 ClassMetaTable.scala 88:49 ClassMetaTable.scala 72:42]
  assign meta_table_io_data_in_a_field_type_4_is_host = _T & io_class_meta_init_bits_desc_state_field_type_4_is_host; // @[ClassMetaTable.scala 85:36 ClassMetaTable.scala 88:49 ClassMetaTable.scala 72:42]
  assign meta_table_io_data_in_a_field_type_5_is_repeated = _T &
    io_class_meta_init_bits_desc_state_field_type_5_is_repeated; // @[ClassMetaTable.scala 85:36 ClassMetaTable.scala 88:49 ClassMetaTable.scala 72:42]
  assign meta_table_io_data_in_a_field_type_5_field_type = _T ?
    io_class_meta_init_bits_desc_state_field_type_5_field_type : 5'h0; // @[ClassMetaTable.scala 85:36 ClassMetaTable.scala 88:49 ClassMetaTable.scala 72:42]
  assign meta_table_io_data_in_a_field_type_5_sub_class_id = _T ?
    io_class_meta_init_bits_desc_state_field_type_5_sub_class_id : 16'h0; // @[ClassMetaTable.scala 85:36 ClassMetaTable.scala 88:49 ClassMetaTable.scala 72:42]
  assign meta_table_io_data_in_a_field_type_5_is_host = _T & io_class_meta_init_bits_desc_state_field_type_5_is_host; // @[ClassMetaTable.scala 85:36 ClassMetaTable.scala 88:49 ClassMetaTable.scala 72:42]
  assign meta_table_io_data_in_a_field_type_6_is_repeated = _T &
    io_class_meta_init_bits_desc_state_field_type_6_is_repeated; // @[ClassMetaTable.scala 85:36 ClassMetaTable.scala 88:49 ClassMetaTable.scala 72:42]
  assign meta_table_io_data_in_a_field_type_6_field_type = _T ?
    io_class_meta_init_bits_desc_state_field_type_6_field_type : 5'h0; // @[ClassMetaTable.scala 85:36 ClassMetaTable.scala 88:49 ClassMetaTable.scala 72:42]
  assign meta_table_io_data_in_a_field_type_6_sub_class_id = _T ?
    io_class_meta_init_bits_desc_state_field_type_6_sub_class_id : 16'h0; // @[ClassMetaTable.scala 85:36 ClassMetaTable.scala 88:49 ClassMetaTable.scala 72:42]
  assign meta_table_io_data_in_a_field_type_6_is_host = _T & io_class_meta_init_bits_desc_state_field_type_6_is_host; // @[ClassMetaTable.scala 85:36 ClassMetaTable.scala 88:49 ClassMetaTable.scala 72:42]
  assign meta_table_io_data_in_a_field_type_7_is_repeated = _T &
    io_class_meta_init_bits_desc_state_field_type_7_is_repeated; // @[ClassMetaTable.scala 85:36 ClassMetaTable.scala 88:49 ClassMetaTable.scala 72:42]
  assign meta_table_io_data_in_a_field_type_7_field_type = _T ?
    io_class_meta_init_bits_desc_state_field_type_7_field_type : 5'h0; // @[ClassMetaTable.scala 85:36 ClassMetaTable.scala 88:49 ClassMetaTable.scala 72:42]
  assign meta_table_io_data_in_a_field_type_7_sub_class_id = _T ?
    io_class_meta_init_bits_desc_state_field_type_7_sub_class_id : 16'h0; // @[ClassMetaTable.scala 85:36 ClassMetaTable.scala 88:49 ClassMetaTable.scala 72:42]
  assign meta_table_io_data_in_a_field_type_7_is_host = _T & io_class_meta_init_bits_desc_state_field_type_7_is_host; // @[ClassMetaTable.scala 85:36 ClassMetaTable.scala 88:49 ClassMetaTable.scala 72:42]
  assign meta_table_io_data_in_a_field_type_8_is_repeated = _T &
    io_class_meta_init_bits_desc_state_field_type_8_is_repeated; // @[ClassMetaTable.scala 85:36 ClassMetaTable.scala 88:49 ClassMetaTable.scala 72:42]
  assign meta_table_io_data_in_a_field_type_8_field_type = _T ?
    io_class_meta_init_bits_desc_state_field_type_8_field_type : 5'h0; // @[ClassMetaTable.scala 85:36 ClassMetaTable.scala 88:49 ClassMetaTable.scala 72:42]
  assign meta_table_io_data_in_a_field_type_8_sub_class_id = _T ?
    io_class_meta_init_bits_desc_state_field_type_8_sub_class_id : 16'h0; // @[ClassMetaTable.scala 85:36 ClassMetaTable.scala 88:49 ClassMetaTable.scala 72:42]
  assign meta_table_io_data_in_a_field_type_8_is_host = _T & io_class_meta_init_bits_desc_state_field_type_8_is_host; // @[ClassMetaTable.scala 85:36 ClassMetaTable.scala 88:49 ClassMetaTable.scala 72:42]
  assign meta_table_io_data_in_a_field_type_9_is_repeated = _T &
    io_class_meta_init_bits_desc_state_field_type_9_is_repeated; // @[ClassMetaTable.scala 85:36 ClassMetaTable.scala 88:49 ClassMetaTable.scala 72:42]
  assign meta_table_io_data_in_a_field_type_9_field_type = _T ?
    io_class_meta_init_bits_desc_state_field_type_9_field_type : 5'h0; // @[ClassMetaTable.scala 85:36 ClassMetaTable.scala 88:49 ClassMetaTable.scala 72:42]
  assign meta_table_io_data_in_a_field_type_9_sub_class_id = _T ?
    io_class_meta_init_bits_desc_state_field_type_9_sub_class_id : 16'h0; // @[ClassMetaTable.scala 85:36 ClassMetaTable.scala 88:49 ClassMetaTable.scala 72:42]
  assign meta_table_io_data_in_a_field_type_9_is_host = _T & io_class_meta_init_bits_desc_state_field_type_9_is_host; // @[ClassMetaTable.scala 85:36 ClassMetaTable.scala 88:49 ClassMetaTable.scala 72:42]
  assign meta_table_io_data_in_a_field_type_10_is_repeated = _T &
    io_class_meta_init_bits_desc_state_field_type_10_is_repeated; // @[ClassMetaTable.scala 85:36 ClassMetaTable.scala 88:49 ClassMetaTable.scala 72:42]
  assign meta_table_io_data_in_a_field_type_10_field_type = _T ?
    io_class_meta_init_bits_desc_state_field_type_10_field_type : 5'h0; // @[ClassMetaTable.scala 85:36 ClassMetaTable.scala 88:49 ClassMetaTable.scala 72:42]
  assign meta_table_io_data_in_a_field_type_10_sub_class_id = _T ?
    io_class_meta_init_bits_desc_state_field_type_10_sub_class_id : 16'h0; // @[ClassMetaTable.scala 85:36 ClassMetaTable.scala 88:49 ClassMetaTable.scala 72:42]
  assign meta_table_io_data_in_a_field_type_10_is_host = _T & io_class_meta_init_bits_desc_state_field_type_10_is_host; // @[ClassMetaTable.scala 85:36 ClassMetaTable.scala 88:49 ClassMetaTable.scala 72:42]
  assign meta_table_io_data_in_a_field_type_11_is_repeated = _T &
    io_class_meta_init_bits_desc_state_field_type_11_is_repeated; // @[ClassMetaTable.scala 85:36 ClassMetaTable.scala 88:49 ClassMetaTable.scala 72:42]
  assign meta_table_io_data_in_a_field_type_11_field_type = _T ?
    io_class_meta_init_bits_desc_state_field_type_11_field_type : 5'h0; // @[ClassMetaTable.scala 85:36 ClassMetaTable.scala 88:49 ClassMetaTable.scala 72:42]
  assign meta_table_io_data_in_a_field_type_11_sub_class_id = _T ?
    io_class_meta_init_bits_desc_state_field_type_11_sub_class_id : 16'h0; // @[ClassMetaTable.scala 85:36 ClassMetaTable.scala 88:49 ClassMetaTable.scala 72:42]
  assign meta_table_io_data_in_a_field_type_11_is_host = _T & io_class_meta_init_bits_desc_state_field_type_11_is_host; // @[ClassMetaTable.scala 85:36 ClassMetaTable.scala 88:49 ClassMetaTable.scala 72:42]
  assign meta_table_io_data_in_a_field_type_12_is_repeated = _T &
    io_class_meta_init_bits_desc_state_field_type_12_is_repeated; // @[ClassMetaTable.scala 85:36 ClassMetaTable.scala 88:49 ClassMetaTable.scala 72:42]
  assign meta_table_io_data_in_a_field_type_12_field_type = _T ?
    io_class_meta_init_bits_desc_state_field_type_12_field_type : 5'h0; // @[ClassMetaTable.scala 85:36 ClassMetaTable.scala 88:49 ClassMetaTable.scala 72:42]
  assign meta_table_io_data_in_a_field_type_12_sub_class_id = _T ?
    io_class_meta_init_bits_desc_state_field_type_12_sub_class_id : 16'h0; // @[ClassMetaTable.scala 85:36 ClassMetaTable.scala 88:49 ClassMetaTable.scala 72:42]
  assign meta_table_io_data_in_a_field_type_12_is_host = _T & io_class_meta_init_bits_desc_state_field_type_12_is_host; // @[ClassMetaTable.scala 85:36 ClassMetaTable.scala 88:49 ClassMetaTable.scala 72:42]
  assign meta_table_io_data_in_a_field_type_13_is_repeated = _T &
    io_class_meta_init_bits_desc_state_field_type_13_is_repeated; // @[ClassMetaTable.scala 85:36 ClassMetaTable.scala 88:49 ClassMetaTable.scala 72:42]
  assign meta_table_io_data_in_a_field_type_13_field_type = _T ?
    io_class_meta_init_bits_desc_state_field_type_13_field_type : 5'h0; // @[ClassMetaTable.scala 85:36 ClassMetaTable.scala 88:49 ClassMetaTable.scala 72:42]
  assign meta_table_io_data_in_a_field_type_13_sub_class_id = _T ?
    io_class_meta_init_bits_desc_state_field_type_13_sub_class_id : 16'h0; // @[ClassMetaTable.scala 85:36 ClassMetaTable.scala 88:49 ClassMetaTable.scala 72:42]
  assign meta_table_io_data_in_a_field_type_13_is_host = _T & io_class_meta_init_bits_desc_state_field_type_13_is_host; // @[ClassMetaTable.scala 85:36 ClassMetaTable.scala 88:49 ClassMetaTable.scala 72:42]
  assign meta_table_io_data_in_a_field_type_14_is_repeated = _T &
    io_class_meta_init_bits_desc_state_field_type_14_is_repeated; // @[ClassMetaTable.scala 85:36 ClassMetaTable.scala 88:49 ClassMetaTable.scala 72:42]
  assign meta_table_io_data_in_a_field_type_14_field_type = _T ?
    io_class_meta_init_bits_desc_state_field_type_14_field_type : 5'h0; // @[ClassMetaTable.scala 85:36 ClassMetaTable.scala 88:49 ClassMetaTable.scala 72:42]
  assign meta_table_io_data_in_a_field_type_14_sub_class_id = _T ?
    io_class_meta_init_bits_desc_state_field_type_14_sub_class_id : 16'h0; // @[ClassMetaTable.scala 85:36 ClassMetaTable.scala 88:49 ClassMetaTable.scala 72:42]
  assign meta_table_io_data_in_a_field_type_14_is_host = _T & io_class_meta_init_bits_desc_state_field_type_14_is_host; // @[ClassMetaTable.scala 85:36 ClassMetaTable.scala 88:49 ClassMetaTable.scala 72:42]
  assign meta_table_io_data_in_a_field_type_15_is_repeated = _T &
    io_class_meta_init_bits_desc_state_field_type_15_is_repeated; // @[ClassMetaTable.scala 85:36 ClassMetaTable.scala 88:49 ClassMetaTable.scala 72:42]
  assign meta_table_io_data_in_a_field_type_15_field_type = _T ?
    io_class_meta_init_bits_desc_state_field_type_15_field_type : 5'h0; // @[ClassMetaTable.scala 85:36 ClassMetaTable.scala 88:49 ClassMetaTable.scala 72:42]
  assign meta_table_io_data_in_a_field_type_15_sub_class_id = _T ?
    io_class_meta_init_bits_desc_state_field_type_15_sub_class_id : 16'h0; // @[ClassMetaTable.scala 85:36 ClassMetaTable.scala 88:49 ClassMetaTable.scala 72:42]
  assign meta_table_io_data_in_a_field_type_15_is_host = _T & io_class_meta_init_bits_desc_state_field_type_15_is_host; // @[ClassMetaTable.scala 85:36 ClassMetaTable.scala 88:49 ClassMetaTable.scala 72:42]
  assign meta_table_io_data_in_a_field_type_16_is_repeated = _T &
    io_class_meta_init_bits_desc_state_field_type_16_is_repeated; // @[ClassMetaTable.scala 85:36 ClassMetaTable.scala 88:49 ClassMetaTable.scala 72:42]
  assign meta_table_io_data_in_a_field_type_16_field_type = _T ?
    io_class_meta_init_bits_desc_state_field_type_16_field_type : 5'h0; // @[ClassMetaTable.scala 85:36 ClassMetaTable.scala 88:49 ClassMetaTable.scala 72:42]
  assign meta_table_io_data_in_a_field_type_16_sub_class_id = _T ?
    io_class_meta_init_bits_desc_state_field_type_16_sub_class_id : 16'h0; // @[ClassMetaTable.scala 85:36 ClassMetaTable.scala 88:49 ClassMetaTable.scala 72:42]
  assign meta_table_io_data_in_a_field_type_16_is_host = _T & io_class_meta_init_bits_desc_state_field_type_16_is_host; // @[ClassMetaTable.scala 85:36 ClassMetaTable.scala 88:49 ClassMetaTable.scala 72:42]
  assign meta_table_io_data_in_a_field_type_17_is_repeated = _T &
    io_class_meta_init_bits_desc_state_field_type_17_is_repeated; // @[ClassMetaTable.scala 85:36 ClassMetaTable.scala 88:49 ClassMetaTable.scala 72:42]
  assign meta_table_io_data_in_a_field_type_17_field_type = _T ?
    io_class_meta_init_bits_desc_state_field_type_17_field_type : 5'h0; // @[ClassMetaTable.scala 85:36 ClassMetaTable.scala 88:49 ClassMetaTable.scala 72:42]
  assign meta_table_io_data_in_a_field_type_17_sub_class_id = _T ?
    io_class_meta_init_bits_desc_state_field_type_17_sub_class_id : 16'h0; // @[ClassMetaTable.scala 85:36 ClassMetaTable.scala 88:49 ClassMetaTable.scala 72:42]
  assign meta_table_io_data_in_a_field_type_17_is_host = _T & io_class_meta_init_bits_desc_state_field_type_17_is_host; // @[ClassMetaTable.scala 85:36 ClassMetaTable.scala 88:49 ClassMetaTable.scala 72:42]
  assign meta_table_io_data_in_a_field_type_18_is_repeated = _T &
    io_class_meta_init_bits_desc_state_field_type_18_is_repeated; // @[ClassMetaTable.scala 85:36 ClassMetaTable.scala 88:49 ClassMetaTable.scala 72:42]
  assign meta_table_io_data_in_a_field_type_18_field_type = _T ?
    io_class_meta_init_bits_desc_state_field_type_18_field_type : 5'h0; // @[ClassMetaTable.scala 85:36 ClassMetaTable.scala 88:49 ClassMetaTable.scala 72:42]
  assign meta_table_io_data_in_a_field_type_18_sub_class_id = _T ?
    io_class_meta_init_bits_desc_state_field_type_18_sub_class_id : 16'h0; // @[ClassMetaTable.scala 85:36 ClassMetaTable.scala 88:49 ClassMetaTable.scala 72:42]
  assign meta_table_io_data_in_a_field_type_18_is_host = _T & io_class_meta_init_bits_desc_state_field_type_18_is_host; // @[ClassMetaTable.scala 85:36 ClassMetaTable.scala 88:49 ClassMetaTable.scala 72:42]
  assign meta_table_io_data_in_a_field_type_19_is_repeated = _T &
    io_class_meta_init_bits_desc_state_field_type_19_is_repeated; // @[ClassMetaTable.scala 85:36 ClassMetaTable.scala 88:49 ClassMetaTable.scala 72:42]
  assign meta_table_io_data_in_a_field_type_19_field_type = _T ?
    io_class_meta_init_bits_desc_state_field_type_19_field_type : 5'h0; // @[ClassMetaTable.scala 85:36 ClassMetaTable.scala 88:49 ClassMetaTable.scala 72:42]
  assign meta_table_io_data_in_a_field_type_19_sub_class_id = _T ?
    io_class_meta_init_bits_desc_state_field_type_19_sub_class_id : 16'h0; // @[ClassMetaTable.scala 85:36 ClassMetaTable.scala 88:49 ClassMetaTable.scala 72:42]
  assign meta_table_io_data_in_a_field_type_19_is_host = _T & io_class_meta_init_bits_desc_state_field_type_19_is_host; // @[ClassMetaTable.scala 85:36 ClassMetaTable.scala 88:49 ClassMetaTable.scala 72:42]
  assign meta_table_io_data_in_a_field_type_20_is_repeated = _T &
    io_class_meta_init_bits_desc_state_field_type_20_is_repeated; // @[ClassMetaTable.scala 85:36 ClassMetaTable.scala 88:49 ClassMetaTable.scala 72:42]
  assign meta_table_io_data_in_a_field_type_20_field_type = _T ?
    io_class_meta_init_bits_desc_state_field_type_20_field_type : 5'h0; // @[ClassMetaTable.scala 85:36 ClassMetaTable.scala 88:49 ClassMetaTable.scala 72:42]
  assign meta_table_io_data_in_a_field_type_20_sub_class_id = _T ?
    io_class_meta_init_bits_desc_state_field_type_20_sub_class_id : 16'h0; // @[ClassMetaTable.scala 85:36 ClassMetaTable.scala 88:49 ClassMetaTable.scala 72:42]
  assign meta_table_io_data_in_a_field_type_20_is_host = _T & io_class_meta_init_bits_desc_state_field_type_20_is_host; // @[ClassMetaTable.scala 85:36 ClassMetaTable.scala 88:49 ClassMetaTable.scala 72:42]
  assign meta_table_io_data_in_a_field_type_21_is_repeated = _T &
    io_class_meta_init_bits_desc_state_field_type_21_is_repeated; // @[ClassMetaTable.scala 85:36 ClassMetaTable.scala 88:49 ClassMetaTable.scala 72:42]
  assign meta_table_io_data_in_a_field_type_21_field_type = _T ?
    io_class_meta_init_bits_desc_state_field_type_21_field_type : 5'h0; // @[ClassMetaTable.scala 85:36 ClassMetaTable.scala 88:49 ClassMetaTable.scala 72:42]
  assign meta_table_io_data_in_a_field_type_21_sub_class_id = _T ?
    io_class_meta_init_bits_desc_state_field_type_21_sub_class_id : 16'h0; // @[ClassMetaTable.scala 85:36 ClassMetaTable.scala 88:49 ClassMetaTable.scala 72:42]
  assign meta_table_io_data_in_a_field_type_21_is_host = _T & io_class_meta_init_bits_desc_state_field_type_21_is_host; // @[ClassMetaTable.scala 85:36 ClassMetaTable.scala 88:49 ClassMetaTable.scala 72:42]
  assign meta_table_io_data_in_a_field_type_22_is_repeated = _T &
    io_class_meta_init_bits_desc_state_field_type_22_is_repeated; // @[ClassMetaTable.scala 85:36 ClassMetaTable.scala 88:49 ClassMetaTable.scala 72:42]
  assign meta_table_io_data_in_a_field_type_22_field_type = _T ?
    io_class_meta_init_bits_desc_state_field_type_22_field_type : 5'h0; // @[ClassMetaTable.scala 85:36 ClassMetaTable.scala 88:49 ClassMetaTable.scala 72:42]
  assign meta_table_io_data_in_a_field_type_22_sub_class_id = _T ?
    io_class_meta_init_bits_desc_state_field_type_22_sub_class_id : 16'h0; // @[ClassMetaTable.scala 85:36 ClassMetaTable.scala 88:49 ClassMetaTable.scala 72:42]
  assign meta_table_io_data_in_a_field_type_22_is_host = _T & io_class_meta_init_bits_desc_state_field_type_22_is_host; // @[ClassMetaTable.scala 85:36 ClassMetaTable.scala 88:49 ClassMetaTable.scala 72:42]
  assign meta_table_io_data_in_a_field_type_23_is_repeated = _T &
    io_class_meta_init_bits_desc_state_field_type_23_is_repeated; // @[ClassMetaTable.scala 85:36 ClassMetaTable.scala 88:49 ClassMetaTable.scala 72:42]
  assign meta_table_io_data_in_a_field_type_23_field_type = _T ?
    io_class_meta_init_bits_desc_state_field_type_23_field_type : 5'h0; // @[ClassMetaTable.scala 85:36 ClassMetaTable.scala 88:49 ClassMetaTable.scala 72:42]
  assign meta_table_io_data_in_a_field_type_23_sub_class_id = _T ?
    io_class_meta_init_bits_desc_state_field_type_23_sub_class_id : 16'h0; // @[ClassMetaTable.scala 85:36 ClassMetaTable.scala 88:49 ClassMetaTable.scala 72:42]
  assign meta_table_io_data_in_a_field_type_23_is_host = _T & io_class_meta_init_bits_desc_state_field_type_23_is_host; // @[ClassMetaTable.scala 85:36 ClassMetaTable.scala 88:49 ClassMetaTable.scala 72:42]
  assign meta_table_io_data_in_a_field_type_24_is_repeated = _T &
    io_class_meta_init_bits_desc_state_field_type_24_is_repeated; // @[ClassMetaTable.scala 85:36 ClassMetaTable.scala 88:49 ClassMetaTable.scala 72:42]
  assign meta_table_io_data_in_a_field_type_24_field_type = _T ?
    io_class_meta_init_bits_desc_state_field_type_24_field_type : 5'h0; // @[ClassMetaTable.scala 85:36 ClassMetaTable.scala 88:49 ClassMetaTable.scala 72:42]
  assign meta_table_io_data_in_a_field_type_24_sub_class_id = _T ?
    io_class_meta_init_bits_desc_state_field_type_24_sub_class_id : 16'h0; // @[ClassMetaTable.scala 85:36 ClassMetaTable.scala 88:49 ClassMetaTable.scala 72:42]
  assign meta_table_io_data_in_a_field_type_24_is_host = _T & io_class_meta_init_bits_desc_state_field_type_24_is_host; // @[ClassMetaTable.scala 85:36 ClassMetaTable.scala 88:49 ClassMetaTable.scala 72:42]
  assign meta_table_io_data_in_a_field_type_25_is_repeated = _T &
    io_class_meta_init_bits_desc_state_field_type_25_is_repeated; // @[ClassMetaTable.scala 85:36 ClassMetaTable.scala 88:49 ClassMetaTable.scala 72:42]
  assign meta_table_io_data_in_a_field_type_25_field_type = _T ?
    io_class_meta_init_bits_desc_state_field_type_25_field_type : 5'h0; // @[ClassMetaTable.scala 85:36 ClassMetaTable.scala 88:49 ClassMetaTable.scala 72:42]
  assign meta_table_io_data_in_a_field_type_25_sub_class_id = _T ?
    io_class_meta_init_bits_desc_state_field_type_25_sub_class_id : 16'h0; // @[ClassMetaTable.scala 85:36 ClassMetaTable.scala 88:49 ClassMetaTable.scala 72:42]
  assign meta_table_io_data_in_a_field_type_25_is_host = _T & io_class_meta_init_bits_desc_state_field_type_25_is_host; // @[ClassMetaTable.scala 85:36 ClassMetaTable.scala 88:49 ClassMetaTable.scala 72:42]
  assign meta_table_io_data_in_a_field_type_26_is_repeated = _T &
    io_class_meta_init_bits_desc_state_field_type_26_is_repeated; // @[ClassMetaTable.scala 85:36 ClassMetaTable.scala 88:49 ClassMetaTable.scala 72:42]
  assign meta_table_io_data_in_a_field_type_26_field_type = _T ?
    io_class_meta_init_bits_desc_state_field_type_26_field_type : 5'h0; // @[ClassMetaTable.scala 85:36 ClassMetaTable.scala 88:49 ClassMetaTable.scala 72:42]
  assign meta_table_io_data_in_a_field_type_26_sub_class_id = _T ?
    io_class_meta_init_bits_desc_state_field_type_26_sub_class_id : 16'h0; // @[ClassMetaTable.scala 85:36 ClassMetaTable.scala 88:49 ClassMetaTable.scala 72:42]
  assign meta_table_io_data_in_a_field_type_26_is_host = _T & io_class_meta_init_bits_desc_state_field_type_26_is_host; // @[ClassMetaTable.scala 85:36 ClassMetaTable.scala 88:49 ClassMetaTable.scala 72:42]
  assign meta_table_io_data_in_a_field_type_27_is_repeated = _T &
    io_class_meta_init_bits_desc_state_field_type_27_is_repeated; // @[ClassMetaTable.scala 85:36 ClassMetaTable.scala 88:49 ClassMetaTable.scala 72:42]
  assign meta_table_io_data_in_a_field_type_27_field_type = _T ?
    io_class_meta_init_bits_desc_state_field_type_27_field_type : 5'h0; // @[ClassMetaTable.scala 85:36 ClassMetaTable.scala 88:49 ClassMetaTable.scala 72:42]
  assign meta_table_io_data_in_a_field_type_27_sub_class_id = _T ?
    io_class_meta_init_bits_desc_state_field_type_27_sub_class_id : 16'h0; // @[ClassMetaTable.scala 85:36 ClassMetaTable.scala 88:49 ClassMetaTable.scala 72:42]
  assign meta_table_io_data_in_a_field_type_27_is_host = _T & io_class_meta_init_bits_desc_state_field_type_27_is_host; // @[ClassMetaTable.scala 85:36 ClassMetaTable.scala 88:49 ClassMetaTable.scala 72:42]
  assign meta_table_io_data_in_a_field_type_28_is_repeated = _T &
    io_class_meta_init_bits_desc_state_field_type_28_is_repeated; // @[ClassMetaTable.scala 85:36 ClassMetaTable.scala 88:49 ClassMetaTable.scala 72:42]
  assign meta_table_io_data_in_a_field_type_28_field_type = _T ?
    io_class_meta_init_bits_desc_state_field_type_28_field_type : 5'h0; // @[ClassMetaTable.scala 85:36 ClassMetaTable.scala 88:49 ClassMetaTable.scala 72:42]
  assign meta_table_io_data_in_a_field_type_28_sub_class_id = _T ?
    io_class_meta_init_bits_desc_state_field_type_28_sub_class_id : 16'h0; // @[ClassMetaTable.scala 85:36 ClassMetaTable.scala 88:49 ClassMetaTable.scala 72:42]
  assign meta_table_io_data_in_a_field_type_28_is_host = _T & io_class_meta_init_bits_desc_state_field_type_28_is_host; // @[ClassMetaTable.scala 85:36 ClassMetaTable.scala 88:49 ClassMetaTable.scala 72:42]
  assign meta_table_io_data_in_a_field_type_29_is_repeated = _T &
    io_class_meta_init_bits_desc_state_field_type_29_is_repeated; // @[ClassMetaTable.scala 85:36 ClassMetaTable.scala 88:49 ClassMetaTable.scala 72:42]
  assign meta_table_io_data_in_a_field_type_29_field_type = _T ?
    io_class_meta_init_bits_desc_state_field_type_29_field_type : 5'h0; // @[ClassMetaTable.scala 85:36 ClassMetaTable.scala 88:49 ClassMetaTable.scala 72:42]
  assign meta_table_io_data_in_a_field_type_29_sub_class_id = _T ?
    io_class_meta_init_bits_desc_state_field_type_29_sub_class_id : 16'h0; // @[ClassMetaTable.scala 85:36 ClassMetaTable.scala 88:49 ClassMetaTable.scala 72:42]
  assign meta_table_io_data_in_a_field_type_29_is_host = _T & io_class_meta_init_bits_desc_state_field_type_29_is_host; // @[ClassMetaTable.scala 85:36 ClassMetaTable.scala 88:49 ClassMetaTable.scala 72:42]
  assign meta_table_io_data_in_a_field_type_30_is_repeated = _T &
    io_class_meta_init_bits_desc_state_field_type_30_is_repeated; // @[ClassMetaTable.scala 85:36 ClassMetaTable.scala 88:49 ClassMetaTable.scala 72:42]
  assign meta_table_io_data_in_a_field_type_30_field_type = _T ?
    io_class_meta_init_bits_desc_state_field_type_30_field_type : 5'h0; // @[ClassMetaTable.scala 85:36 ClassMetaTable.scala 88:49 ClassMetaTable.scala 72:42]
  assign meta_table_io_data_in_a_field_type_30_sub_class_id = _T ?
    io_class_meta_init_bits_desc_state_field_type_30_sub_class_id : 16'h0; // @[ClassMetaTable.scala 85:36 ClassMetaTable.scala 88:49 ClassMetaTable.scala 72:42]
  assign meta_table_io_data_in_a_field_type_30_is_host = _T & io_class_meta_init_bits_desc_state_field_type_30_is_host; // @[ClassMetaTable.scala 85:36 ClassMetaTable.scala 88:49 ClassMetaTable.scala 72:42]
  assign meta_table_io_data_in_a_field_type_31_is_repeated = _T &
    io_class_meta_init_bits_desc_state_field_type_31_is_repeated; // @[ClassMetaTable.scala 85:36 ClassMetaTable.scala 88:49 ClassMetaTable.scala 72:42]
  assign meta_table_io_data_in_a_field_type_31_field_type = _T ?
    io_class_meta_init_bits_desc_state_field_type_31_field_type : 5'h0; // @[ClassMetaTable.scala 85:36 ClassMetaTable.scala 88:49 ClassMetaTable.scala 72:42]
  assign meta_table_io_data_in_a_field_type_31_sub_class_id = _T ?
    io_class_meta_init_bits_desc_state_field_type_31_sub_class_id : 16'h0; // @[ClassMetaTable.scala 85:36 ClassMetaTable.scala 88:49 ClassMetaTable.scala 72:42]
  assign meta_table_io_data_in_a_field_type_31_is_host = _T & io_class_meta_init_bits_desc_state_field_type_31_is_host; // @[ClassMetaTable.scala 85:36 ClassMetaTable.scala 88:49 ClassMetaTable.scala 72:42]
  assign meta_table_io_data_in_a_field_type_32_is_repeated = _T &
    io_class_meta_init_bits_desc_state_field_type_32_is_repeated; // @[ClassMetaTable.scala 85:36 ClassMetaTable.scala 88:49 ClassMetaTable.scala 72:42]
  assign meta_table_io_data_in_a_field_type_32_field_type = _T ?
    io_class_meta_init_bits_desc_state_field_type_32_field_type : 5'h0; // @[ClassMetaTable.scala 85:36 ClassMetaTable.scala 88:49 ClassMetaTable.scala 72:42]
  assign meta_table_io_data_in_a_field_type_32_sub_class_id = _T ?
    io_class_meta_init_bits_desc_state_field_type_32_sub_class_id : 16'h0; // @[ClassMetaTable.scala 85:36 ClassMetaTable.scala 88:49 ClassMetaTable.scala 72:42]
  assign meta_table_io_data_in_a_field_type_32_is_host = _T & io_class_meta_init_bits_desc_state_field_type_32_is_host; // @[ClassMetaTable.scala 85:36 ClassMetaTable.scala 88:49 ClassMetaTable.scala 72:42]
  always @(posedge clock) begin
    if (reset) begin // @[Collector.scala 169:42]
      counter <= 32'h0; // @[Collector.scala 169:42]
    end else if (_T) begin // @[Collector.scala 170:34]
      counter <= _counter_T_1; // @[Collector.scala 171:41]
    end
    if (reset) begin // @[ClassMetaTable.scala 67:46]
      state <= 2'h0; // @[ClassMetaTable.scala 67:46]
    end else if (_T) begin // @[ClassMetaTable.scala 85:36]
      state <= 2'h0; // @[ClassMetaTable.scala 89:49]
    end else if (_T_2) begin // @[ClassMetaTable.scala 90:52]
      state <= 2'h1; // @[ClassMetaTable.scala 93:49]
    end else if (_T_3) begin // @[ClassMetaTable.scala 94:52]
      state <= 2'h2; // @[ClassMetaTable.scala 97:49]
    end else begin
      state <= 2'h0; // @[ClassMetaTable.scala 99:49]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  counter = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  state = _RAND_1[1:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Control(
  input          clock,
  input          reset,
  output         io_axi_aw_ready,
  input          io_axi_aw_valid,
  input  [63:0]  io_axi_aw_bits_addr,
  output         io_axi_w_ready,
  input          io_axi_w_valid,
  input  [511:0] io_axi_w_bits_data,
  input          io_axi_r_ready,
  output         io_axi_r_valid,
  output [511:0] io_axi_r_bits_data,
  output         io_metadata_init_valid,
  output [9:0]   io_metadata_init_bits_class_id,
  output [15:0]  io_metadata_init_bits_desc_state_class_length,
  output [7:0]   io_metadata_init_bits_desc_state_max_field_num,
  output         io_metadata_init_bits_desc_state_field_type_0_is_repeated,
  output [4:0]   io_metadata_init_bits_desc_state_field_type_0_field_type,
  output [15:0]  io_metadata_init_bits_desc_state_field_type_0_sub_class_id,
  output         io_metadata_init_bits_desc_state_field_type_0_is_host,
  output         io_metadata_init_bits_desc_state_field_type_1_is_repeated,
  output [4:0]   io_metadata_init_bits_desc_state_field_type_1_field_type,
  output [15:0]  io_metadata_init_bits_desc_state_field_type_1_sub_class_id,
  output         io_metadata_init_bits_desc_state_field_type_1_is_host,
  output         io_metadata_init_bits_desc_state_field_type_2_is_repeated,
  output [4:0]   io_metadata_init_bits_desc_state_field_type_2_field_type,
  output [15:0]  io_metadata_init_bits_desc_state_field_type_2_sub_class_id,
  output         io_metadata_init_bits_desc_state_field_type_2_is_host,
  output         io_metadata_init_bits_desc_state_field_type_3_is_repeated,
  output [4:0]   io_metadata_init_bits_desc_state_field_type_3_field_type,
  output [15:0]  io_metadata_init_bits_desc_state_field_type_3_sub_class_id,
  output         io_metadata_init_bits_desc_state_field_type_3_is_host,
  output         io_metadata_init_bits_desc_state_field_type_4_is_repeated,
  output [4:0]   io_metadata_init_bits_desc_state_field_type_4_field_type,
  output [15:0]  io_metadata_init_bits_desc_state_field_type_4_sub_class_id,
  output         io_metadata_init_bits_desc_state_field_type_4_is_host,
  output         io_metadata_init_bits_desc_state_field_type_5_is_repeated,
  output [4:0]   io_metadata_init_bits_desc_state_field_type_5_field_type,
  output [15:0]  io_metadata_init_bits_desc_state_field_type_5_sub_class_id,
  output         io_metadata_init_bits_desc_state_field_type_5_is_host,
  output         io_metadata_init_bits_desc_state_field_type_6_is_repeated,
  output [4:0]   io_metadata_init_bits_desc_state_field_type_6_field_type,
  output [15:0]  io_metadata_init_bits_desc_state_field_type_6_sub_class_id,
  output         io_metadata_init_bits_desc_state_field_type_6_is_host,
  output         io_metadata_init_bits_desc_state_field_type_7_is_repeated,
  output [4:0]   io_metadata_init_bits_desc_state_field_type_7_field_type,
  output [15:0]  io_metadata_init_bits_desc_state_field_type_7_sub_class_id,
  output         io_metadata_init_bits_desc_state_field_type_7_is_host,
  output         io_metadata_init_bits_desc_state_field_type_8_is_repeated,
  output [4:0]   io_metadata_init_bits_desc_state_field_type_8_field_type,
  output [15:0]  io_metadata_init_bits_desc_state_field_type_8_sub_class_id,
  output         io_metadata_init_bits_desc_state_field_type_8_is_host,
  output         io_metadata_init_bits_desc_state_field_type_9_is_repeated,
  output [4:0]   io_metadata_init_bits_desc_state_field_type_9_field_type,
  output [15:0]  io_metadata_init_bits_desc_state_field_type_9_sub_class_id,
  output         io_metadata_init_bits_desc_state_field_type_9_is_host,
  output         io_metadata_init_bits_desc_state_field_type_10_is_repeated,
  output [4:0]   io_metadata_init_bits_desc_state_field_type_10_field_type,
  output [15:0]  io_metadata_init_bits_desc_state_field_type_10_sub_class_id,
  output         io_metadata_init_bits_desc_state_field_type_10_is_host,
  output         io_metadata_init_bits_desc_state_field_type_11_is_repeated,
  output [4:0]   io_metadata_init_bits_desc_state_field_type_11_field_type,
  output [15:0]  io_metadata_init_bits_desc_state_field_type_11_sub_class_id,
  output         io_metadata_init_bits_desc_state_field_type_11_is_host,
  output         io_metadata_init_bits_desc_state_field_type_12_is_repeated,
  output [4:0]   io_metadata_init_bits_desc_state_field_type_12_field_type,
  output [15:0]  io_metadata_init_bits_desc_state_field_type_12_sub_class_id,
  output         io_metadata_init_bits_desc_state_field_type_12_is_host,
  output         io_metadata_init_bits_desc_state_field_type_13_is_repeated,
  output [4:0]   io_metadata_init_bits_desc_state_field_type_13_field_type,
  output [15:0]  io_metadata_init_bits_desc_state_field_type_13_sub_class_id,
  output         io_metadata_init_bits_desc_state_field_type_13_is_host,
  output         io_metadata_init_bits_desc_state_field_type_14_is_repeated,
  output [4:0]   io_metadata_init_bits_desc_state_field_type_14_field_type,
  output [15:0]  io_metadata_init_bits_desc_state_field_type_14_sub_class_id,
  output         io_metadata_init_bits_desc_state_field_type_14_is_host,
  output         io_metadata_init_bits_desc_state_field_type_15_is_repeated,
  output [4:0]   io_metadata_init_bits_desc_state_field_type_15_field_type,
  output [15:0]  io_metadata_init_bits_desc_state_field_type_15_sub_class_id,
  output         io_metadata_init_bits_desc_state_field_type_15_is_host,
  output         io_metadata_init_bits_desc_state_field_type_16_is_repeated,
  output [4:0]   io_metadata_init_bits_desc_state_field_type_16_field_type,
  output [15:0]  io_metadata_init_bits_desc_state_field_type_16_sub_class_id,
  output         io_metadata_init_bits_desc_state_field_type_16_is_host,
  output         io_metadata_init_bits_desc_state_field_type_17_is_repeated,
  output [4:0]   io_metadata_init_bits_desc_state_field_type_17_field_type,
  output [15:0]  io_metadata_init_bits_desc_state_field_type_17_sub_class_id,
  output         io_metadata_init_bits_desc_state_field_type_17_is_host,
  output         io_metadata_init_bits_desc_state_field_type_18_is_repeated,
  output [4:0]   io_metadata_init_bits_desc_state_field_type_18_field_type,
  output [15:0]  io_metadata_init_bits_desc_state_field_type_18_sub_class_id,
  output         io_metadata_init_bits_desc_state_field_type_18_is_host,
  output         io_metadata_init_bits_desc_state_field_type_19_is_repeated,
  output [4:0]   io_metadata_init_bits_desc_state_field_type_19_field_type,
  output [15:0]  io_metadata_init_bits_desc_state_field_type_19_sub_class_id,
  output         io_metadata_init_bits_desc_state_field_type_19_is_host,
  output         io_metadata_init_bits_desc_state_field_type_20_is_repeated,
  output [4:0]   io_metadata_init_bits_desc_state_field_type_20_field_type,
  output [15:0]  io_metadata_init_bits_desc_state_field_type_20_sub_class_id,
  output         io_metadata_init_bits_desc_state_field_type_20_is_host,
  output         io_metadata_init_bits_desc_state_field_type_21_is_repeated,
  output [4:0]   io_metadata_init_bits_desc_state_field_type_21_field_type,
  output [15:0]  io_metadata_init_bits_desc_state_field_type_21_sub_class_id,
  output         io_metadata_init_bits_desc_state_field_type_21_is_host,
  output         io_metadata_init_bits_desc_state_field_type_22_is_repeated,
  output [4:0]   io_metadata_init_bits_desc_state_field_type_22_field_type,
  output [15:0]  io_metadata_init_bits_desc_state_field_type_22_sub_class_id,
  output         io_metadata_init_bits_desc_state_field_type_22_is_host,
  output         io_metadata_init_bits_desc_state_field_type_23_is_repeated,
  output [4:0]   io_metadata_init_bits_desc_state_field_type_23_field_type,
  output [15:0]  io_metadata_init_bits_desc_state_field_type_23_sub_class_id,
  output         io_metadata_init_bits_desc_state_field_type_23_is_host,
  output         io_metadata_init_bits_desc_state_field_type_24_is_repeated,
  output [4:0]   io_metadata_init_bits_desc_state_field_type_24_field_type,
  output [15:0]  io_metadata_init_bits_desc_state_field_type_24_sub_class_id,
  output         io_metadata_init_bits_desc_state_field_type_24_is_host,
  output         io_metadata_init_bits_desc_state_field_type_25_is_repeated,
  output [4:0]   io_metadata_init_bits_desc_state_field_type_25_field_type,
  output [15:0]  io_metadata_init_bits_desc_state_field_type_25_sub_class_id,
  output         io_metadata_init_bits_desc_state_field_type_25_is_host,
  output         io_metadata_init_bits_desc_state_field_type_26_is_repeated,
  output [4:0]   io_metadata_init_bits_desc_state_field_type_26_field_type,
  output [15:0]  io_metadata_init_bits_desc_state_field_type_26_sub_class_id,
  output         io_metadata_init_bits_desc_state_field_type_26_is_host,
  output         io_metadata_init_bits_desc_state_field_type_27_is_repeated,
  output [4:0]   io_metadata_init_bits_desc_state_field_type_27_field_type,
  output [15:0]  io_metadata_init_bits_desc_state_field_type_27_sub_class_id,
  output         io_metadata_init_bits_desc_state_field_type_27_is_host,
  output         io_metadata_init_bits_desc_state_field_type_28_is_repeated,
  output [4:0]   io_metadata_init_bits_desc_state_field_type_28_field_type,
  output [15:0]  io_metadata_init_bits_desc_state_field_type_28_sub_class_id,
  output         io_metadata_init_bits_desc_state_field_type_28_is_host,
  output         io_metadata_init_bits_desc_state_field_type_29_is_repeated,
  output [4:0]   io_metadata_init_bits_desc_state_field_type_29_field_type,
  output [15:0]  io_metadata_init_bits_desc_state_field_type_29_sub_class_id,
  output         io_metadata_init_bits_desc_state_field_type_29_is_host,
  output         io_metadata_init_bits_desc_state_field_type_30_is_repeated,
  output [4:0]   io_metadata_init_bits_desc_state_field_type_30_field_type,
  output [15:0]  io_metadata_init_bits_desc_state_field_type_30_sub_class_id,
  output         io_metadata_init_bits_desc_state_field_type_30_is_host,
  output         io_metadata_init_bits_desc_state_field_type_31_is_repeated,
  output [4:0]   io_metadata_init_bits_desc_state_field_type_31_field_type,
  output [15:0]  io_metadata_init_bits_desc_state_field_type_31_sub_class_id,
  output         io_metadata_init_bits_desc_state_field_type_31_is_host,
  output         io_metadata_init_bits_desc_state_field_type_32_is_repeated,
  output [4:0]   io_metadata_init_bits_desc_state_field_type_32_field_type,
  output [15:0]  io_metadata_init_bits_desc_state_field_type_32_sub_class_id,
  output         io_metadata_init_bits_desc_state_field_type_32_is_host,
  input          io_ser_cmd_ready,
  output         io_ser_cmd_valid,
  output [9:0]   io_ser_cmd_bits_class_id,
  output [63:0]  io_ser_cmd_bits_host_base_addr
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
`endif // RANDOMIZE_REG_INIT
  reg [2:0] s_wr; // @[Control.scala 43:27]
  reg [31:0] cur_data; // @[Control.scala 56:31]
  reg [9:0] classmeta_reg_class_id; // @[Control.scala 57:36]
  reg [15:0] classmeta_reg_desc_state_class_length; // @[Control.scala 57:36]
  reg [7:0] classmeta_reg_desc_state_max_field_num; // @[Control.scala 57:36]
  reg  classmeta_reg_desc_state_field_type_0_is_repeated; // @[Control.scala 57:36]
  reg [4:0] classmeta_reg_desc_state_field_type_0_field_type; // @[Control.scala 57:36]
  reg [15:0] classmeta_reg_desc_state_field_type_0_sub_class_id; // @[Control.scala 57:36]
  reg  classmeta_reg_desc_state_field_type_0_is_host; // @[Control.scala 57:36]
  reg  classmeta_reg_desc_state_field_type_1_is_repeated; // @[Control.scala 57:36]
  reg [4:0] classmeta_reg_desc_state_field_type_1_field_type; // @[Control.scala 57:36]
  reg [15:0] classmeta_reg_desc_state_field_type_1_sub_class_id; // @[Control.scala 57:36]
  reg  classmeta_reg_desc_state_field_type_1_is_host; // @[Control.scala 57:36]
  reg  classmeta_reg_desc_state_field_type_2_is_repeated; // @[Control.scala 57:36]
  reg [4:0] classmeta_reg_desc_state_field_type_2_field_type; // @[Control.scala 57:36]
  reg [15:0] classmeta_reg_desc_state_field_type_2_sub_class_id; // @[Control.scala 57:36]
  reg  classmeta_reg_desc_state_field_type_2_is_host; // @[Control.scala 57:36]
  reg  classmeta_reg_desc_state_field_type_3_is_repeated; // @[Control.scala 57:36]
  reg [4:0] classmeta_reg_desc_state_field_type_3_field_type; // @[Control.scala 57:36]
  reg [15:0] classmeta_reg_desc_state_field_type_3_sub_class_id; // @[Control.scala 57:36]
  reg  classmeta_reg_desc_state_field_type_3_is_host; // @[Control.scala 57:36]
  reg  classmeta_reg_desc_state_field_type_4_is_repeated; // @[Control.scala 57:36]
  reg [4:0] classmeta_reg_desc_state_field_type_4_field_type; // @[Control.scala 57:36]
  reg [15:0] classmeta_reg_desc_state_field_type_4_sub_class_id; // @[Control.scala 57:36]
  reg  classmeta_reg_desc_state_field_type_4_is_host; // @[Control.scala 57:36]
  reg  classmeta_reg_desc_state_field_type_5_is_repeated; // @[Control.scala 57:36]
  reg [4:0] classmeta_reg_desc_state_field_type_5_field_type; // @[Control.scala 57:36]
  reg [15:0] classmeta_reg_desc_state_field_type_5_sub_class_id; // @[Control.scala 57:36]
  reg  classmeta_reg_desc_state_field_type_5_is_host; // @[Control.scala 57:36]
  reg  classmeta_reg_desc_state_field_type_6_is_repeated; // @[Control.scala 57:36]
  reg [4:0] classmeta_reg_desc_state_field_type_6_field_type; // @[Control.scala 57:36]
  reg [15:0] classmeta_reg_desc_state_field_type_6_sub_class_id; // @[Control.scala 57:36]
  reg  classmeta_reg_desc_state_field_type_6_is_host; // @[Control.scala 57:36]
  reg  classmeta_reg_desc_state_field_type_7_is_repeated; // @[Control.scala 57:36]
  reg [4:0] classmeta_reg_desc_state_field_type_7_field_type; // @[Control.scala 57:36]
  reg [15:0] classmeta_reg_desc_state_field_type_7_sub_class_id; // @[Control.scala 57:36]
  reg  classmeta_reg_desc_state_field_type_7_is_host; // @[Control.scala 57:36]
  reg  classmeta_reg_desc_state_field_type_8_is_repeated; // @[Control.scala 57:36]
  reg [4:0] classmeta_reg_desc_state_field_type_8_field_type; // @[Control.scala 57:36]
  reg [15:0] classmeta_reg_desc_state_field_type_8_sub_class_id; // @[Control.scala 57:36]
  reg  classmeta_reg_desc_state_field_type_8_is_host; // @[Control.scala 57:36]
  reg  classmeta_reg_desc_state_field_type_9_is_repeated; // @[Control.scala 57:36]
  reg [4:0] classmeta_reg_desc_state_field_type_9_field_type; // @[Control.scala 57:36]
  reg [15:0] classmeta_reg_desc_state_field_type_9_sub_class_id; // @[Control.scala 57:36]
  reg  classmeta_reg_desc_state_field_type_9_is_host; // @[Control.scala 57:36]
  reg  classmeta_reg_desc_state_field_type_10_is_repeated; // @[Control.scala 57:36]
  reg [4:0] classmeta_reg_desc_state_field_type_10_field_type; // @[Control.scala 57:36]
  reg [15:0] classmeta_reg_desc_state_field_type_10_sub_class_id; // @[Control.scala 57:36]
  reg  classmeta_reg_desc_state_field_type_10_is_host; // @[Control.scala 57:36]
  reg  classmeta_reg_desc_state_field_type_11_is_repeated; // @[Control.scala 57:36]
  reg [4:0] classmeta_reg_desc_state_field_type_11_field_type; // @[Control.scala 57:36]
  reg [15:0] classmeta_reg_desc_state_field_type_11_sub_class_id; // @[Control.scala 57:36]
  reg  classmeta_reg_desc_state_field_type_11_is_host; // @[Control.scala 57:36]
  reg  classmeta_reg_desc_state_field_type_12_is_repeated; // @[Control.scala 57:36]
  reg [4:0] classmeta_reg_desc_state_field_type_12_field_type; // @[Control.scala 57:36]
  reg [15:0] classmeta_reg_desc_state_field_type_12_sub_class_id; // @[Control.scala 57:36]
  reg  classmeta_reg_desc_state_field_type_12_is_host; // @[Control.scala 57:36]
  reg  classmeta_reg_desc_state_field_type_13_is_repeated; // @[Control.scala 57:36]
  reg [4:0] classmeta_reg_desc_state_field_type_13_field_type; // @[Control.scala 57:36]
  reg [15:0] classmeta_reg_desc_state_field_type_13_sub_class_id; // @[Control.scala 57:36]
  reg  classmeta_reg_desc_state_field_type_13_is_host; // @[Control.scala 57:36]
  reg  classmeta_reg_desc_state_field_type_14_is_repeated; // @[Control.scala 57:36]
  reg [4:0] classmeta_reg_desc_state_field_type_14_field_type; // @[Control.scala 57:36]
  reg [15:0] classmeta_reg_desc_state_field_type_14_sub_class_id; // @[Control.scala 57:36]
  reg  classmeta_reg_desc_state_field_type_14_is_host; // @[Control.scala 57:36]
  reg  classmeta_reg_desc_state_field_type_15_is_repeated; // @[Control.scala 57:36]
  reg [4:0] classmeta_reg_desc_state_field_type_15_field_type; // @[Control.scala 57:36]
  reg [15:0] classmeta_reg_desc_state_field_type_15_sub_class_id; // @[Control.scala 57:36]
  reg  classmeta_reg_desc_state_field_type_15_is_host; // @[Control.scala 57:36]
  reg  classmeta_reg_desc_state_field_type_16_is_repeated; // @[Control.scala 57:36]
  reg [4:0] classmeta_reg_desc_state_field_type_16_field_type; // @[Control.scala 57:36]
  reg [15:0] classmeta_reg_desc_state_field_type_16_sub_class_id; // @[Control.scala 57:36]
  reg  classmeta_reg_desc_state_field_type_16_is_host; // @[Control.scala 57:36]
  reg  classmeta_reg_desc_state_field_type_17_is_repeated; // @[Control.scala 57:36]
  reg [4:0] classmeta_reg_desc_state_field_type_17_field_type; // @[Control.scala 57:36]
  reg [15:0] classmeta_reg_desc_state_field_type_17_sub_class_id; // @[Control.scala 57:36]
  reg  classmeta_reg_desc_state_field_type_17_is_host; // @[Control.scala 57:36]
  reg  classmeta_reg_desc_state_field_type_18_is_repeated; // @[Control.scala 57:36]
  reg [4:0] classmeta_reg_desc_state_field_type_18_field_type; // @[Control.scala 57:36]
  reg [15:0] classmeta_reg_desc_state_field_type_18_sub_class_id; // @[Control.scala 57:36]
  reg  classmeta_reg_desc_state_field_type_18_is_host; // @[Control.scala 57:36]
  reg  classmeta_reg_desc_state_field_type_19_is_repeated; // @[Control.scala 57:36]
  reg [4:0] classmeta_reg_desc_state_field_type_19_field_type; // @[Control.scala 57:36]
  reg [15:0] classmeta_reg_desc_state_field_type_19_sub_class_id; // @[Control.scala 57:36]
  reg  classmeta_reg_desc_state_field_type_19_is_host; // @[Control.scala 57:36]
  reg  classmeta_reg_desc_state_field_type_20_is_repeated; // @[Control.scala 57:36]
  reg [4:0] classmeta_reg_desc_state_field_type_20_field_type; // @[Control.scala 57:36]
  reg [15:0] classmeta_reg_desc_state_field_type_20_sub_class_id; // @[Control.scala 57:36]
  reg  classmeta_reg_desc_state_field_type_20_is_host; // @[Control.scala 57:36]
  reg  classmeta_reg_desc_state_field_type_21_is_repeated; // @[Control.scala 57:36]
  reg [4:0] classmeta_reg_desc_state_field_type_21_field_type; // @[Control.scala 57:36]
  reg [15:0] classmeta_reg_desc_state_field_type_21_sub_class_id; // @[Control.scala 57:36]
  reg  classmeta_reg_desc_state_field_type_21_is_host; // @[Control.scala 57:36]
  reg  classmeta_reg_desc_state_field_type_22_is_repeated; // @[Control.scala 57:36]
  reg [4:0] classmeta_reg_desc_state_field_type_22_field_type; // @[Control.scala 57:36]
  reg [15:0] classmeta_reg_desc_state_field_type_22_sub_class_id; // @[Control.scala 57:36]
  reg  classmeta_reg_desc_state_field_type_22_is_host; // @[Control.scala 57:36]
  reg  classmeta_reg_desc_state_field_type_23_is_repeated; // @[Control.scala 57:36]
  reg [4:0] classmeta_reg_desc_state_field_type_23_field_type; // @[Control.scala 57:36]
  reg [15:0] classmeta_reg_desc_state_field_type_23_sub_class_id; // @[Control.scala 57:36]
  reg  classmeta_reg_desc_state_field_type_23_is_host; // @[Control.scala 57:36]
  reg  classmeta_reg_desc_state_field_type_24_is_repeated; // @[Control.scala 57:36]
  reg [4:0] classmeta_reg_desc_state_field_type_24_field_type; // @[Control.scala 57:36]
  reg [15:0] classmeta_reg_desc_state_field_type_24_sub_class_id; // @[Control.scala 57:36]
  reg  classmeta_reg_desc_state_field_type_24_is_host; // @[Control.scala 57:36]
  reg  classmeta_reg_desc_state_field_type_25_is_repeated; // @[Control.scala 57:36]
  reg [4:0] classmeta_reg_desc_state_field_type_25_field_type; // @[Control.scala 57:36]
  reg [15:0] classmeta_reg_desc_state_field_type_25_sub_class_id; // @[Control.scala 57:36]
  reg  classmeta_reg_desc_state_field_type_25_is_host; // @[Control.scala 57:36]
  reg  classmeta_reg_desc_state_field_type_26_is_repeated; // @[Control.scala 57:36]
  reg [4:0] classmeta_reg_desc_state_field_type_26_field_type; // @[Control.scala 57:36]
  reg [15:0] classmeta_reg_desc_state_field_type_26_sub_class_id; // @[Control.scala 57:36]
  reg  classmeta_reg_desc_state_field_type_26_is_host; // @[Control.scala 57:36]
  reg  classmeta_reg_desc_state_field_type_27_is_repeated; // @[Control.scala 57:36]
  reg [4:0] classmeta_reg_desc_state_field_type_27_field_type; // @[Control.scala 57:36]
  reg [15:0] classmeta_reg_desc_state_field_type_27_sub_class_id; // @[Control.scala 57:36]
  reg  classmeta_reg_desc_state_field_type_27_is_host; // @[Control.scala 57:36]
  reg  classmeta_reg_desc_state_field_type_28_is_repeated; // @[Control.scala 57:36]
  reg [4:0] classmeta_reg_desc_state_field_type_28_field_type; // @[Control.scala 57:36]
  reg [15:0] classmeta_reg_desc_state_field_type_28_sub_class_id; // @[Control.scala 57:36]
  reg  classmeta_reg_desc_state_field_type_28_is_host; // @[Control.scala 57:36]
  reg  classmeta_reg_desc_state_field_type_29_is_repeated; // @[Control.scala 57:36]
  reg [4:0] classmeta_reg_desc_state_field_type_29_field_type; // @[Control.scala 57:36]
  reg [15:0] classmeta_reg_desc_state_field_type_29_sub_class_id; // @[Control.scala 57:36]
  reg  classmeta_reg_desc_state_field_type_29_is_host; // @[Control.scala 57:36]
  wire  _T = io_axi_r_ready & io_axi_r_valid; // @[Decoupled.scala 40:37]
  wire [31:0] _cur_data_T_1 = cur_data + 32'h1; // @[Control.scala 59:38]
  wire  _T_1 = 3'h0 == s_wr; // @[Conditional.scala 37:30]
  wire  _T_2 = io_axi_aw_ready & io_axi_aw_valid; // @[Decoupled.scala 40:37]
  wire [63:0] _w_addr_T = {{6'd0}, io_axi_aw_bits_addr[63:6]}; // @[Control.scala 75:73]
  wire [2:0] _GEN_1 = _w_addr_T == 64'hd ? 3'h7 : 3'h1; // @[Control.scala 86:84 Control.scala 87:53 Control.scala 89:33]
  wire [2:0] _GEN_2 = _w_addr_T == 64'hc ? 3'h6 : _GEN_1; // @[Control.scala 84:84 Control.scala 85:53]
  wire [2:0] _GEN_3 = _w_addr_T == 64'h16 ? 3'h5 : _GEN_2; // @[Control.scala 82:87 Control.scala 83:53]
  wire [2:0] _GEN_4 = _w_addr_T == 64'h15 ? 3'h4 : _GEN_3; // @[Control.scala 80:87 Control.scala 81:53]
  wire [2:0] _GEN_5 = _w_addr_T == 64'h14 ? 3'h3 : _GEN_4; // @[Control.scala 78:71 Control.scala 79:53]
  wire  _T_15 = 3'h2 == s_wr; // @[Conditional.scala 37:30]
  wire  _T_16 = io_axi_w_ready & io_axi_w_valid; // @[Decoupled.scala 40:37]
  wire [2:0] _GEN_11 = _T_16 ? 3'h0 : s_wr; // @[Control.scala 94:39 Control.scala 97:57 Control.scala 43:27]
  wire  _T_17 = 3'h3 == s_wr; // @[Conditional.scala 37:30]
  wire [10:0] _GEN_12 = _T_16 ? io_axi_w_bits_data[10:0] : {{1'd0}, classmeta_reg_class_id}; // @[Control.scala 101:39 Control.scala 102:45 Control.scala 57:36]
  wire [15:0] _GEN_13 = _T_16 ? io_axi_w_bits_data[31:16] : {{8'd0}, classmeta_reg_desc_state_max_field_num}; // @[Control.scala 101:39 Control.scala 103:56 Control.scala 57:36]
  wire [31:0] _GEN_14 = _T_16 ? io_axi_w_bits_data[63:32] : {{16'd0}, classmeta_reg_desc_state_class_length}; // @[Control.scala 101:39 Control.scala 104:73 Control.scala 57:36]
  wire  _GEN_15 = _T_16 ? io_axi_w_bits_data[64] : classmeta_reg_desc_state_field_type_0_is_host; // @[Control.scala 101:39 Control.scala 106:75 Control.scala 57:36]
  wire  _GEN_16 = _T_16 ? io_axi_w_bits_data[65] : classmeta_reg_desc_state_field_type_0_is_repeated; // @[Control.scala 101:39 Control.scala 107:75 Control.scala 57:36]
  wire [4:0] _GEN_17 = _T_16 ? io_axi_w_bits_data[70:66] : classmeta_reg_desc_state_field_type_0_field_type; // @[Control.scala 101:39 Control.scala 108:75 Control.scala 57:36]
  wire [15:0] _GEN_18 = _T_16 ? io_axi_w_bits_data[95:80] : classmeta_reg_desc_state_field_type_0_sub_class_id; // @[Control.scala 101:39 Control.scala 109:75 Control.scala 57:36]
  wire  _GEN_19 = _T_16 ? io_axi_w_bits_data[96] : classmeta_reg_desc_state_field_type_1_is_host; // @[Control.scala 101:39 Control.scala 106:75 Control.scala 57:36]
  wire  _GEN_20 = _T_16 ? io_axi_w_bits_data[97] : classmeta_reg_desc_state_field_type_1_is_repeated; // @[Control.scala 101:39 Control.scala 107:75 Control.scala 57:36]
  wire [4:0] _GEN_21 = _T_16 ? io_axi_w_bits_data[102:98] : classmeta_reg_desc_state_field_type_1_field_type; // @[Control.scala 101:39 Control.scala 108:75 Control.scala 57:36]
  wire [15:0] _GEN_22 = _T_16 ? io_axi_w_bits_data[127:112] : classmeta_reg_desc_state_field_type_1_sub_class_id; // @[Control.scala 101:39 Control.scala 109:75 Control.scala 57:36]
  wire  _GEN_23 = _T_16 ? io_axi_w_bits_data[128] : classmeta_reg_desc_state_field_type_2_is_host; // @[Control.scala 101:39 Control.scala 106:75 Control.scala 57:36]
  wire  _GEN_24 = _T_16 ? io_axi_w_bits_data[129] : classmeta_reg_desc_state_field_type_2_is_repeated; // @[Control.scala 101:39 Control.scala 107:75 Control.scala 57:36]
  wire [4:0] _GEN_25 = _T_16 ? io_axi_w_bits_data[134:130] : classmeta_reg_desc_state_field_type_2_field_type; // @[Control.scala 101:39 Control.scala 108:75 Control.scala 57:36]
  wire [15:0] _GEN_26 = _T_16 ? io_axi_w_bits_data[159:144] : classmeta_reg_desc_state_field_type_2_sub_class_id; // @[Control.scala 101:39 Control.scala 109:75 Control.scala 57:36]
  wire  _GEN_27 = _T_16 ? io_axi_w_bits_data[160] : classmeta_reg_desc_state_field_type_3_is_host; // @[Control.scala 101:39 Control.scala 106:75 Control.scala 57:36]
  wire  _GEN_28 = _T_16 ? io_axi_w_bits_data[161] : classmeta_reg_desc_state_field_type_3_is_repeated; // @[Control.scala 101:39 Control.scala 107:75 Control.scala 57:36]
  wire [4:0] _GEN_29 = _T_16 ? io_axi_w_bits_data[166:162] : classmeta_reg_desc_state_field_type_3_field_type; // @[Control.scala 101:39 Control.scala 108:75 Control.scala 57:36]
  wire [15:0] _GEN_30 = _T_16 ? io_axi_w_bits_data[191:176] : classmeta_reg_desc_state_field_type_3_sub_class_id; // @[Control.scala 101:39 Control.scala 109:75 Control.scala 57:36]
  wire  _GEN_31 = _T_16 ? io_axi_w_bits_data[192] : classmeta_reg_desc_state_field_type_4_is_host; // @[Control.scala 101:39 Control.scala 106:75 Control.scala 57:36]
  wire  _GEN_32 = _T_16 ? io_axi_w_bits_data[193] : classmeta_reg_desc_state_field_type_4_is_repeated; // @[Control.scala 101:39 Control.scala 107:75 Control.scala 57:36]
  wire [4:0] _GEN_33 = _T_16 ? io_axi_w_bits_data[198:194] : classmeta_reg_desc_state_field_type_4_field_type; // @[Control.scala 101:39 Control.scala 108:75 Control.scala 57:36]
  wire [15:0] _GEN_34 = _T_16 ? io_axi_w_bits_data[223:208] : classmeta_reg_desc_state_field_type_4_sub_class_id; // @[Control.scala 101:39 Control.scala 109:75 Control.scala 57:36]
  wire  _GEN_35 = _T_16 ? io_axi_w_bits_data[224] : classmeta_reg_desc_state_field_type_5_is_host; // @[Control.scala 101:39 Control.scala 106:75 Control.scala 57:36]
  wire  _GEN_36 = _T_16 ? io_axi_w_bits_data[225] : classmeta_reg_desc_state_field_type_5_is_repeated; // @[Control.scala 101:39 Control.scala 107:75 Control.scala 57:36]
  wire [4:0] _GEN_37 = _T_16 ? io_axi_w_bits_data[230:226] : classmeta_reg_desc_state_field_type_5_field_type; // @[Control.scala 101:39 Control.scala 108:75 Control.scala 57:36]
  wire [15:0] _GEN_38 = _T_16 ? io_axi_w_bits_data[255:240] : classmeta_reg_desc_state_field_type_5_sub_class_id; // @[Control.scala 101:39 Control.scala 109:75 Control.scala 57:36]
  wire  _GEN_39 = _T_16 ? io_axi_w_bits_data[256] : classmeta_reg_desc_state_field_type_6_is_host; // @[Control.scala 101:39 Control.scala 106:75 Control.scala 57:36]
  wire  _GEN_40 = _T_16 ? io_axi_w_bits_data[257] : classmeta_reg_desc_state_field_type_6_is_repeated; // @[Control.scala 101:39 Control.scala 107:75 Control.scala 57:36]
  wire [4:0] _GEN_41 = _T_16 ? io_axi_w_bits_data[262:258] : classmeta_reg_desc_state_field_type_6_field_type; // @[Control.scala 101:39 Control.scala 108:75 Control.scala 57:36]
  wire [15:0] _GEN_42 = _T_16 ? io_axi_w_bits_data[287:272] : classmeta_reg_desc_state_field_type_6_sub_class_id; // @[Control.scala 101:39 Control.scala 109:75 Control.scala 57:36]
  wire  _GEN_43 = _T_16 ? io_axi_w_bits_data[288] : classmeta_reg_desc_state_field_type_7_is_host; // @[Control.scala 101:39 Control.scala 106:75 Control.scala 57:36]
  wire  _GEN_44 = _T_16 ? io_axi_w_bits_data[289] : classmeta_reg_desc_state_field_type_7_is_repeated; // @[Control.scala 101:39 Control.scala 107:75 Control.scala 57:36]
  wire [4:0] _GEN_45 = _T_16 ? io_axi_w_bits_data[294:290] : classmeta_reg_desc_state_field_type_7_field_type; // @[Control.scala 101:39 Control.scala 108:75 Control.scala 57:36]
  wire [15:0] _GEN_46 = _T_16 ? io_axi_w_bits_data[319:304] : classmeta_reg_desc_state_field_type_7_sub_class_id; // @[Control.scala 101:39 Control.scala 109:75 Control.scala 57:36]
  wire  _GEN_47 = _T_16 ? io_axi_w_bits_data[320] : classmeta_reg_desc_state_field_type_8_is_host; // @[Control.scala 101:39 Control.scala 106:75 Control.scala 57:36]
  wire  _GEN_48 = _T_16 ? io_axi_w_bits_data[321] : classmeta_reg_desc_state_field_type_8_is_repeated; // @[Control.scala 101:39 Control.scala 107:75 Control.scala 57:36]
  wire [4:0] _GEN_49 = _T_16 ? io_axi_w_bits_data[326:322] : classmeta_reg_desc_state_field_type_8_field_type; // @[Control.scala 101:39 Control.scala 108:75 Control.scala 57:36]
  wire [15:0] _GEN_50 = _T_16 ? io_axi_w_bits_data[351:336] : classmeta_reg_desc_state_field_type_8_sub_class_id; // @[Control.scala 101:39 Control.scala 109:75 Control.scala 57:36]
  wire  _GEN_51 = _T_16 ? io_axi_w_bits_data[352] : classmeta_reg_desc_state_field_type_9_is_host; // @[Control.scala 101:39 Control.scala 106:75 Control.scala 57:36]
  wire  _GEN_52 = _T_16 ? io_axi_w_bits_data[353] : classmeta_reg_desc_state_field_type_9_is_repeated; // @[Control.scala 101:39 Control.scala 107:75 Control.scala 57:36]
  wire [4:0] _GEN_53 = _T_16 ? io_axi_w_bits_data[358:354] : classmeta_reg_desc_state_field_type_9_field_type; // @[Control.scala 101:39 Control.scala 108:75 Control.scala 57:36]
  wire [15:0] _GEN_54 = _T_16 ? io_axi_w_bits_data[383:368] : classmeta_reg_desc_state_field_type_9_sub_class_id; // @[Control.scala 101:39 Control.scala 109:75 Control.scala 57:36]
  wire  _GEN_55 = _T_16 ? io_axi_w_bits_data[384] : classmeta_reg_desc_state_field_type_10_is_host; // @[Control.scala 101:39 Control.scala 106:75 Control.scala 57:36]
  wire  _GEN_56 = _T_16 ? io_axi_w_bits_data[385] : classmeta_reg_desc_state_field_type_10_is_repeated; // @[Control.scala 101:39 Control.scala 107:75 Control.scala 57:36]
  wire [4:0] _GEN_57 = _T_16 ? io_axi_w_bits_data[390:386] : classmeta_reg_desc_state_field_type_10_field_type; // @[Control.scala 101:39 Control.scala 108:75 Control.scala 57:36]
  wire [15:0] _GEN_58 = _T_16 ? io_axi_w_bits_data[415:400] : classmeta_reg_desc_state_field_type_10_sub_class_id; // @[Control.scala 101:39 Control.scala 109:75 Control.scala 57:36]
  wire  _GEN_59 = _T_16 ? io_axi_w_bits_data[416] : classmeta_reg_desc_state_field_type_11_is_host; // @[Control.scala 101:39 Control.scala 106:75 Control.scala 57:36]
  wire  _GEN_60 = _T_16 ? io_axi_w_bits_data[417] : classmeta_reg_desc_state_field_type_11_is_repeated; // @[Control.scala 101:39 Control.scala 107:75 Control.scala 57:36]
  wire [4:0] _GEN_61 = _T_16 ? io_axi_w_bits_data[422:418] : classmeta_reg_desc_state_field_type_11_field_type; // @[Control.scala 101:39 Control.scala 108:75 Control.scala 57:36]
  wire [15:0] _GEN_62 = _T_16 ? io_axi_w_bits_data[447:432] : classmeta_reg_desc_state_field_type_11_sub_class_id; // @[Control.scala 101:39 Control.scala 109:75 Control.scala 57:36]
  wire  _GEN_63 = _T_16 ? io_axi_w_bits_data[448] : classmeta_reg_desc_state_field_type_12_is_host; // @[Control.scala 101:39 Control.scala 106:75 Control.scala 57:36]
  wire  _GEN_64 = _T_16 ? io_axi_w_bits_data[449] : classmeta_reg_desc_state_field_type_12_is_repeated; // @[Control.scala 101:39 Control.scala 107:75 Control.scala 57:36]
  wire [4:0] _GEN_65 = _T_16 ? io_axi_w_bits_data[454:450] : classmeta_reg_desc_state_field_type_12_field_type; // @[Control.scala 101:39 Control.scala 108:75 Control.scala 57:36]
  wire [15:0] _GEN_66 = _T_16 ? io_axi_w_bits_data[479:464] : classmeta_reg_desc_state_field_type_12_sub_class_id; // @[Control.scala 101:39 Control.scala 109:75 Control.scala 57:36]
  wire  _GEN_67 = _T_16 ? io_axi_w_bits_data[480] : classmeta_reg_desc_state_field_type_13_is_host; // @[Control.scala 101:39 Control.scala 106:75 Control.scala 57:36]
  wire  _GEN_68 = _T_16 ? io_axi_w_bits_data[481] : classmeta_reg_desc_state_field_type_13_is_repeated; // @[Control.scala 101:39 Control.scala 107:75 Control.scala 57:36]
  wire [4:0] _GEN_69 = _T_16 ? io_axi_w_bits_data[486:482] : classmeta_reg_desc_state_field_type_13_field_type; // @[Control.scala 101:39 Control.scala 108:75 Control.scala 57:36]
  wire [15:0] _GEN_70 = _T_16 ? io_axi_w_bits_data[511:496] : classmeta_reg_desc_state_field_type_13_sub_class_id; // @[Control.scala 101:39 Control.scala 109:75 Control.scala 57:36]
  wire  _T_19 = 3'h4 == s_wr; // @[Conditional.scala 37:30]
  wire  _GEN_72 = _T_16 ? io_axi_w_bits_data[0] : classmeta_reg_desc_state_field_type_14_is_host; // @[Control.scala 115:39 Control.scala 117:76 Control.scala 57:36]
  wire  _GEN_73 = _T_16 ? io_axi_w_bits_data[1] : classmeta_reg_desc_state_field_type_14_is_repeated; // @[Control.scala 115:39 Control.scala 118:76 Control.scala 57:36]
  wire [4:0] _GEN_74 = _T_16 ? io_axi_w_bits_data[6:2] : classmeta_reg_desc_state_field_type_14_field_type; // @[Control.scala 115:39 Control.scala 119:76 Control.scala 57:36]
  wire [15:0] _GEN_75 = _T_16 ? io_axi_w_bits_data[31:16] : classmeta_reg_desc_state_field_type_14_sub_class_id; // @[Control.scala 115:39 Control.scala 120:76 Control.scala 57:36]
  wire  _GEN_76 = _T_16 ? io_axi_w_bits_data[32] : classmeta_reg_desc_state_field_type_15_is_host; // @[Control.scala 115:39 Control.scala 117:76 Control.scala 57:36]
  wire  _GEN_77 = _T_16 ? io_axi_w_bits_data[33] : classmeta_reg_desc_state_field_type_15_is_repeated; // @[Control.scala 115:39 Control.scala 118:76 Control.scala 57:36]
  wire [4:0] _GEN_78 = _T_16 ? io_axi_w_bits_data[38:34] : classmeta_reg_desc_state_field_type_15_field_type; // @[Control.scala 115:39 Control.scala 119:76 Control.scala 57:36]
  wire [15:0] _GEN_79 = _T_16 ? io_axi_w_bits_data[63:48] : classmeta_reg_desc_state_field_type_15_sub_class_id; // @[Control.scala 115:39 Control.scala 120:76 Control.scala 57:36]
  wire  _GEN_80 = _T_16 ? io_axi_w_bits_data[64] : classmeta_reg_desc_state_field_type_16_is_host; // @[Control.scala 115:39 Control.scala 117:76 Control.scala 57:36]
  wire  _GEN_81 = _T_16 ? io_axi_w_bits_data[65] : classmeta_reg_desc_state_field_type_16_is_repeated; // @[Control.scala 115:39 Control.scala 118:76 Control.scala 57:36]
  wire [4:0] _GEN_82 = _T_16 ? io_axi_w_bits_data[70:66] : classmeta_reg_desc_state_field_type_16_field_type; // @[Control.scala 115:39 Control.scala 119:76 Control.scala 57:36]
  wire [15:0] _GEN_83 = _T_16 ? io_axi_w_bits_data[95:80] : classmeta_reg_desc_state_field_type_16_sub_class_id; // @[Control.scala 115:39 Control.scala 120:76 Control.scala 57:36]
  wire  _GEN_84 = _T_16 ? io_axi_w_bits_data[96] : classmeta_reg_desc_state_field_type_17_is_host; // @[Control.scala 115:39 Control.scala 117:76 Control.scala 57:36]
  wire  _GEN_85 = _T_16 ? io_axi_w_bits_data[97] : classmeta_reg_desc_state_field_type_17_is_repeated; // @[Control.scala 115:39 Control.scala 118:76 Control.scala 57:36]
  wire [4:0] _GEN_86 = _T_16 ? io_axi_w_bits_data[102:98] : classmeta_reg_desc_state_field_type_17_field_type; // @[Control.scala 115:39 Control.scala 119:76 Control.scala 57:36]
  wire [15:0] _GEN_87 = _T_16 ? io_axi_w_bits_data[127:112] : classmeta_reg_desc_state_field_type_17_sub_class_id; // @[Control.scala 115:39 Control.scala 120:76 Control.scala 57:36]
  wire  _GEN_88 = _T_16 ? io_axi_w_bits_data[128] : classmeta_reg_desc_state_field_type_18_is_host; // @[Control.scala 115:39 Control.scala 117:76 Control.scala 57:36]
  wire  _GEN_89 = _T_16 ? io_axi_w_bits_data[129] : classmeta_reg_desc_state_field_type_18_is_repeated; // @[Control.scala 115:39 Control.scala 118:76 Control.scala 57:36]
  wire [4:0] _GEN_90 = _T_16 ? io_axi_w_bits_data[134:130] : classmeta_reg_desc_state_field_type_18_field_type; // @[Control.scala 115:39 Control.scala 119:76 Control.scala 57:36]
  wire [15:0] _GEN_91 = _T_16 ? io_axi_w_bits_data[159:144] : classmeta_reg_desc_state_field_type_18_sub_class_id; // @[Control.scala 115:39 Control.scala 120:76 Control.scala 57:36]
  wire  _GEN_92 = _T_16 ? io_axi_w_bits_data[160] : classmeta_reg_desc_state_field_type_19_is_host; // @[Control.scala 115:39 Control.scala 117:76 Control.scala 57:36]
  wire  _GEN_93 = _T_16 ? io_axi_w_bits_data[161] : classmeta_reg_desc_state_field_type_19_is_repeated; // @[Control.scala 115:39 Control.scala 118:76 Control.scala 57:36]
  wire [4:0] _GEN_94 = _T_16 ? io_axi_w_bits_data[166:162] : classmeta_reg_desc_state_field_type_19_field_type; // @[Control.scala 115:39 Control.scala 119:76 Control.scala 57:36]
  wire [15:0] _GEN_95 = _T_16 ? io_axi_w_bits_data[191:176] : classmeta_reg_desc_state_field_type_19_sub_class_id; // @[Control.scala 115:39 Control.scala 120:76 Control.scala 57:36]
  wire  _GEN_96 = _T_16 ? io_axi_w_bits_data[192] : classmeta_reg_desc_state_field_type_20_is_host; // @[Control.scala 115:39 Control.scala 117:76 Control.scala 57:36]
  wire  _GEN_97 = _T_16 ? io_axi_w_bits_data[193] : classmeta_reg_desc_state_field_type_20_is_repeated; // @[Control.scala 115:39 Control.scala 118:76 Control.scala 57:36]
  wire [4:0] _GEN_98 = _T_16 ? io_axi_w_bits_data[198:194] : classmeta_reg_desc_state_field_type_20_field_type; // @[Control.scala 115:39 Control.scala 119:76 Control.scala 57:36]
  wire [15:0] _GEN_99 = _T_16 ? io_axi_w_bits_data[223:208] : classmeta_reg_desc_state_field_type_20_sub_class_id; // @[Control.scala 115:39 Control.scala 120:76 Control.scala 57:36]
  wire  _GEN_100 = _T_16 ? io_axi_w_bits_data[224] : classmeta_reg_desc_state_field_type_21_is_host; // @[Control.scala 115:39 Control.scala 117:76 Control.scala 57:36]
  wire  _GEN_101 = _T_16 ? io_axi_w_bits_data[225] : classmeta_reg_desc_state_field_type_21_is_repeated; // @[Control.scala 115:39 Control.scala 118:76 Control.scala 57:36]
  wire [4:0] _GEN_102 = _T_16 ? io_axi_w_bits_data[230:226] : classmeta_reg_desc_state_field_type_21_field_type; // @[Control.scala 115:39 Control.scala 119:76 Control.scala 57:36]
  wire [15:0] _GEN_103 = _T_16 ? io_axi_w_bits_data[255:240] : classmeta_reg_desc_state_field_type_21_sub_class_id; // @[Control.scala 115:39 Control.scala 120:76 Control.scala 57:36]
  wire  _GEN_104 = _T_16 ? io_axi_w_bits_data[256] : classmeta_reg_desc_state_field_type_22_is_host; // @[Control.scala 115:39 Control.scala 117:76 Control.scala 57:36]
  wire  _GEN_105 = _T_16 ? io_axi_w_bits_data[257] : classmeta_reg_desc_state_field_type_22_is_repeated; // @[Control.scala 115:39 Control.scala 118:76 Control.scala 57:36]
  wire [4:0] _GEN_106 = _T_16 ? io_axi_w_bits_data[262:258] : classmeta_reg_desc_state_field_type_22_field_type; // @[Control.scala 115:39 Control.scala 119:76 Control.scala 57:36]
  wire [15:0] _GEN_107 = _T_16 ? io_axi_w_bits_data[287:272] : classmeta_reg_desc_state_field_type_22_sub_class_id; // @[Control.scala 115:39 Control.scala 120:76 Control.scala 57:36]
  wire  _GEN_108 = _T_16 ? io_axi_w_bits_data[288] : classmeta_reg_desc_state_field_type_23_is_host; // @[Control.scala 115:39 Control.scala 117:76 Control.scala 57:36]
  wire  _GEN_109 = _T_16 ? io_axi_w_bits_data[289] : classmeta_reg_desc_state_field_type_23_is_repeated; // @[Control.scala 115:39 Control.scala 118:76 Control.scala 57:36]
  wire [4:0] _GEN_110 = _T_16 ? io_axi_w_bits_data[294:290] : classmeta_reg_desc_state_field_type_23_field_type; // @[Control.scala 115:39 Control.scala 119:76 Control.scala 57:36]
  wire [15:0] _GEN_111 = _T_16 ? io_axi_w_bits_data[319:304] : classmeta_reg_desc_state_field_type_23_sub_class_id; // @[Control.scala 115:39 Control.scala 120:76 Control.scala 57:36]
  wire  _GEN_112 = _T_16 ? io_axi_w_bits_data[320] : classmeta_reg_desc_state_field_type_24_is_host; // @[Control.scala 115:39 Control.scala 117:76 Control.scala 57:36]
  wire  _GEN_113 = _T_16 ? io_axi_w_bits_data[321] : classmeta_reg_desc_state_field_type_24_is_repeated; // @[Control.scala 115:39 Control.scala 118:76 Control.scala 57:36]
  wire [4:0] _GEN_114 = _T_16 ? io_axi_w_bits_data[326:322] : classmeta_reg_desc_state_field_type_24_field_type; // @[Control.scala 115:39 Control.scala 119:76 Control.scala 57:36]
  wire [15:0] _GEN_115 = _T_16 ? io_axi_w_bits_data[351:336] : classmeta_reg_desc_state_field_type_24_sub_class_id; // @[Control.scala 115:39 Control.scala 120:76 Control.scala 57:36]
  wire  _GEN_116 = _T_16 ? io_axi_w_bits_data[352] : classmeta_reg_desc_state_field_type_25_is_host; // @[Control.scala 115:39 Control.scala 117:76 Control.scala 57:36]
  wire  _GEN_117 = _T_16 ? io_axi_w_bits_data[353] : classmeta_reg_desc_state_field_type_25_is_repeated; // @[Control.scala 115:39 Control.scala 118:76 Control.scala 57:36]
  wire [4:0] _GEN_118 = _T_16 ? io_axi_w_bits_data[358:354] : classmeta_reg_desc_state_field_type_25_field_type; // @[Control.scala 115:39 Control.scala 119:76 Control.scala 57:36]
  wire [15:0] _GEN_119 = _T_16 ? io_axi_w_bits_data[383:368] : classmeta_reg_desc_state_field_type_25_sub_class_id; // @[Control.scala 115:39 Control.scala 120:76 Control.scala 57:36]
  wire  _GEN_120 = _T_16 ? io_axi_w_bits_data[384] : classmeta_reg_desc_state_field_type_26_is_host; // @[Control.scala 115:39 Control.scala 117:76 Control.scala 57:36]
  wire  _GEN_121 = _T_16 ? io_axi_w_bits_data[385] : classmeta_reg_desc_state_field_type_26_is_repeated; // @[Control.scala 115:39 Control.scala 118:76 Control.scala 57:36]
  wire [4:0] _GEN_122 = _T_16 ? io_axi_w_bits_data[390:386] : classmeta_reg_desc_state_field_type_26_field_type; // @[Control.scala 115:39 Control.scala 119:76 Control.scala 57:36]
  wire [15:0] _GEN_123 = _T_16 ? io_axi_w_bits_data[415:400] : classmeta_reg_desc_state_field_type_26_sub_class_id; // @[Control.scala 115:39 Control.scala 120:76 Control.scala 57:36]
  wire  _GEN_124 = _T_16 ? io_axi_w_bits_data[416] : classmeta_reg_desc_state_field_type_27_is_host; // @[Control.scala 115:39 Control.scala 117:76 Control.scala 57:36]
  wire  _GEN_125 = _T_16 ? io_axi_w_bits_data[417] : classmeta_reg_desc_state_field_type_27_is_repeated; // @[Control.scala 115:39 Control.scala 118:76 Control.scala 57:36]
  wire [4:0] _GEN_126 = _T_16 ? io_axi_w_bits_data[422:418] : classmeta_reg_desc_state_field_type_27_field_type; // @[Control.scala 115:39 Control.scala 119:76 Control.scala 57:36]
  wire [15:0] _GEN_127 = _T_16 ? io_axi_w_bits_data[447:432] : classmeta_reg_desc_state_field_type_27_sub_class_id; // @[Control.scala 115:39 Control.scala 120:76 Control.scala 57:36]
  wire  _GEN_128 = _T_16 ? io_axi_w_bits_data[448] : classmeta_reg_desc_state_field_type_28_is_host; // @[Control.scala 115:39 Control.scala 117:76 Control.scala 57:36]
  wire  _GEN_129 = _T_16 ? io_axi_w_bits_data[449] : classmeta_reg_desc_state_field_type_28_is_repeated; // @[Control.scala 115:39 Control.scala 118:76 Control.scala 57:36]
  wire [4:0] _GEN_130 = _T_16 ? io_axi_w_bits_data[454:450] : classmeta_reg_desc_state_field_type_28_field_type; // @[Control.scala 115:39 Control.scala 119:76 Control.scala 57:36]
  wire [15:0] _GEN_131 = _T_16 ? io_axi_w_bits_data[479:464] : classmeta_reg_desc_state_field_type_28_sub_class_id; // @[Control.scala 115:39 Control.scala 120:76 Control.scala 57:36]
  wire  _GEN_132 = _T_16 ? io_axi_w_bits_data[480] : classmeta_reg_desc_state_field_type_29_is_host; // @[Control.scala 115:39 Control.scala 117:76 Control.scala 57:36]
  wire  _GEN_133 = _T_16 ? io_axi_w_bits_data[481] : classmeta_reg_desc_state_field_type_29_is_repeated; // @[Control.scala 115:39 Control.scala 118:76 Control.scala 57:36]
  wire [4:0] _GEN_134 = _T_16 ? io_axi_w_bits_data[486:482] : classmeta_reg_desc_state_field_type_29_field_type; // @[Control.scala 115:39 Control.scala 119:76 Control.scala 57:36]
  wire [15:0] _GEN_135 = _T_16 ? io_axi_w_bits_data[511:496] : classmeta_reg_desc_state_field_type_29_sub_class_id; // @[Control.scala 115:39 Control.scala 120:76 Control.scala 57:36]
  wire  _T_21 = 3'h5 == s_wr; // @[Conditional.scala 37:30]
  wire  _GEN_138 = _T_16 & classmeta_reg_desc_state_field_type_0_is_host; // @[Control.scala 126:39 Control.scala 128:65 Util.scala 13:25]
  wire [15:0] _GEN_139 = _T_16 ? classmeta_reg_desc_state_field_type_0_sub_class_id : 16'h0; // @[Control.scala 126:39 Control.scala 128:65 Util.scala 13:25]
  wire [4:0] _GEN_140 = _T_16 ? classmeta_reg_desc_state_field_type_0_field_type : 5'h0; // @[Control.scala 126:39 Control.scala 128:65 Util.scala 13:25]
  wire  _GEN_141 = _T_16 & classmeta_reg_desc_state_field_type_0_is_repeated; // @[Control.scala 126:39 Control.scala 128:65 Util.scala 13:25]
  wire  _GEN_142 = _T_16 & classmeta_reg_desc_state_field_type_1_is_host; // @[Control.scala 126:39 Control.scala 128:65 Util.scala 13:25]
  wire [15:0] _GEN_143 = _T_16 ? classmeta_reg_desc_state_field_type_1_sub_class_id : 16'h0; // @[Control.scala 126:39 Control.scala 128:65 Util.scala 13:25]
  wire [4:0] _GEN_144 = _T_16 ? classmeta_reg_desc_state_field_type_1_field_type : 5'h0; // @[Control.scala 126:39 Control.scala 128:65 Util.scala 13:25]
  wire  _GEN_145 = _T_16 & classmeta_reg_desc_state_field_type_1_is_repeated; // @[Control.scala 126:39 Control.scala 128:65 Util.scala 13:25]
  wire  _GEN_146 = _T_16 & classmeta_reg_desc_state_field_type_2_is_host; // @[Control.scala 126:39 Control.scala 128:65 Util.scala 13:25]
  wire [15:0] _GEN_147 = _T_16 ? classmeta_reg_desc_state_field_type_2_sub_class_id : 16'h0; // @[Control.scala 126:39 Control.scala 128:65 Util.scala 13:25]
  wire [4:0] _GEN_148 = _T_16 ? classmeta_reg_desc_state_field_type_2_field_type : 5'h0; // @[Control.scala 126:39 Control.scala 128:65 Util.scala 13:25]
  wire  _GEN_149 = _T_16 & classmeta_reg_desc_state_field_type_2_is_repeated; // @[Control.scala 126:39 Control.scala 128:65 Util.scala 13:25]
  wire  _GEN_150 = _T_16 & classmeta_reg_desc_state_field_type_3_is_host; // @[Control.scala 126:39 Control.scala 128:65 Util.scala 13:25]
  wire [15:0] _GEN_151 = _T_16 ? classmeta_reg_desc_state_field_type_3_sub_class_id : 16'h0; // @[Control.scala 126:39 Control.scala 128:65 Util.scala 13:25]
  wire [4:0] _GEN_152 = _T_16 ? classmeta_reg_desc_state_field_type_3_field_type : 5'h0; // @[Control.scala 126:39 Control.scala 128:65 Util.scala 13:25]
  wire  _GEN_153 = _T_16 & classmeta_reg_desc_state_field_type_3_is_repeated; // @[Control.scala 126:39 Control.scala 128:65 Util.scala 13:25]
  wire  _GEN_154 = _T_16 & classmeta_reg_desc_state_field_type_4_is_host; // @[Control.scala 126:39 Control.scala 128:65 Util.scala 13:25]
  wire [15:0] _GEN_155 = _T_16 ? classmeta_reg_desc_state_field_type_4_sub_class_id : 16'h0; // @[Control.scala 126:39 Control.scala 128:65 Util.scala 13:25]
  wire [4:0] _GEN_156 = _T_16 ? classmeta_reg_desc_state_field_type_4_field_type : 5'h0; // @[Control.scala 126:39 Control.scala 128:65 Util.scala 13:25]
  wire  _GEN_157 = _T_16 & classmeta_reg_desc_state_field_type_4_is_repeated; // @[Control.scala 126:39 Control.scala 128:65 Util.scala 13:25]
  wire  _GEN_158 = _T_16 & classmeta_reg_desc_state_field_type_5_is_host; // @[Control.scala 126:39 Control.scala 128:65 Util.scala 13:25]
  wire [15:0] _GEN_159 = _T_16 ? classmeta_reg_desc_state_field_type_5_sub_class_id : 16'h0; // @[Control.scala 126:39 Control.scala 128:65 Util.scala 13:25]
  wire [4:0] _GEN_160 = _T_16 ? classmeta_reg_desc_state_field_type_5_field_type : 5'h0; // @[Control.scala 126:39 Control.scala 128:65 Util.scala 13:25]
  wire  _GEN_161 = _T_16 & classmeta_reg_desc_state_field_type_5_is_repeated; // @[Control.scala 126:39 Control.scala 128:65 Util.scala 13:25]
  wire  _GEN_162 = _T_16 & classmeta_reg_desc_state_field_type_6_is_host; // @[Control.scala 126:39 Control.scala 128:65 Util.scala 13:25]
  wire [15:0] _GEN_163 = _T_16 ? classmeta_reg_desc_state_field_type_6_sub_class_id : 16'h0; // @[Control.scala 126:39 Control.scala 128:65 Util.scala 13:25]
  wire [4:0] _GEN_164 = _T_16 ? classmeta_reg_desc_state_field_type_6_field_type : 5'h0; // @[Control.scala 126:39 Control.scala 128:65 Util.scala 13:25]
  wire  _GEN_165 = _T_16 & classmeta_reg_desc_state_field_type_6_is_repeated; // @[Control.scala 126:39 Control.scala 128:65 Util.scala 13:25]
  wire  _GEN_166 = _T_16 & classmeta_reg_desc_state_field_type_7_is_host; // @[Control.scala 126:39 Control.scala 128:65 Util.scala 13:25]
  wire [15:0] _GEN_167 = _T_16 ? classmeta_reg_desc_state_field_type_7_sub_class_id : 16'h0; // @[Control.scala 126:39 Control.scala 128:65 Util.scala 13:25]
  wire [4:0] _GEN_168 = _T_16 ? classmeta_reg_desc_state_field_type_7_field_type : 5'h0; // @[Control.scala 126:39 Control.scala 128:65 Util.scala 13:25]
  wire  _GEN_169 = _T_16 & classmeta_reg_desc_state_field_type_7_is_repeated; // @[Control.scala 126:39 Control.scala 128:65 Util.scala 13:25]
  wire  _GEN_170 = _T_16 & classmeta_reg_desc_state_field_type_8_is_host; // @[Control.scala 126:39 Control.scala 128:65 Util.scala 13:25]
  wire [15:0] _GEN_171 = _T_16 ? classmeta_reg_desc_state_field_type_8_sub_class_id : 16'h0; // @[Control.scala 126:39 Control.scala 128:65 Util.scala 13:25]
  wire [4:0] _GEN_172 = _T_16 ? classmeta_reg_desc_state_field_type_8_field_type : 5'h0; // @[Control.scala 126:39 Control.scala 128:65 Util.scala 13:25]
  wire  _GEN_173 = _T_16 & classmeta_reg_desc_state_field_type_8_is_repeated; // @[Control.scala 126:39 Control.scala 128:65 Util.scala 13:25]
  wire  _GEN_174 = _T_16 & classmeta_reg_desc_state_field_type_9_is_host; // @[Control.scala 126:39 Control.scala 128:65 Util.scala 13:25]
  wire [15:0] _GEN_175 = _T_16 ? classmeta_reg_desc_state_field_type_9_sub_class_id : 16'h0; // @[Control.scala 126:39 Control.scala 128:65 Util.scala 13:25]
  wire [4:0] _GEN_176 = _T_16 ? classmeta_reg_desc_state_field_type_9_field_type : 5'h0; // @[Control.scala 126:39 Control.scala 128:65 Util.scala 13:25]
  wire  _GEN_177 = _T_16 & classmeta_reg_desc_state_field_type_9_is_repeated; // @[Control.scala 126:39 Control.scala 128:65 Util.scala 13:25]
  wire  _GEN_178 = _T_16 & classmeta_reg_desc_state_field_type_10_is_host; // @[Control.scala 126:39 Control.scala 128:65 Util.scala 13:25]
  wire [15:0] _GEN_179 = _T_16 ? classmeta_reg_desc_state_field_type_10_sub_class_id : 16'h0; // @[Control.scala 126:39 Control.scala 128:65 Util.scala 13:25]
  wire [4:0] _GEN_180 = _T_16 ? classmeta_reg_desc_state_field_type_10_field_type : 5'h0; // @[Control.scala 126:39 Control.scala 128:65 Util.scala 13:25]
  wire  _GEN_181 = _T_16 & classmeta_reg_desc_state_field_type_10_is_repeated; // @[Control.scala 126:39 Control.scala 128:65 Util.scala 13:25]
  wire  _GEN_182 = _T_16 & classmeta_reg_desc_state_field_type_11_is_host; // @[Control.scala 126:39 Control.scala 128:65 Util.scala 13:25]
  wire [15:0] _GEN_183 = _T_16 ? classmeta_reg_desc_state_field_type_11_sub_class_id : 16'h0; // @[Control.scala 126:39 Control.scala 128:65 Util.scala 13:25]
  wire [4:0] _GEN_184 = _T_16 ? classmeta_reg_desc_state_field_type_11_field_type : 5'h0; // @[Control.scala 126:39 Control.scala 128:65 Util.scala 13:25]
  wire  _GEN_185 = _T_16 & classmeta_reg_desc_state_field_type_11_is_repeated; // @[Control.scala 126:39 Control.scala 128:65 Util.scala 13:25]
  wire  _GEN_186 = _T_16 & classmeta_reg_desc_state_field_type_12_is_host; // @[Control.scala 126:39 Control.scala 128:65 Util.scala 13:25]
  wire [15:0] _GEN_187 = _T_16 ? classmeta_reg_desc_state_field_type_12_sub_class_id : 16'h0; // @[Control.scala 126:39 Control.scala 128:65 Util.scala 13:25]
  wire [4:0] _GEN_188 = _T_16 ? classmeta_reg_desc_state_field_type_12_field_type : 5'h0; // @[Control.scala 126:39 Control.scala 128:65 Util.scala 13:25]
  wire  _GEN_189 = _T_16 & classmeta_reg_desc_state_field_type_12_is_repeated; // @[Control.scala 126:39 Control.scala 128:65 Util.scala 13:25]
  wire  _GEN_190 = _T_16 & classmeta_reg_desc_state_field_type_13_is_host; // @[Control.scala 126:39 Control.scala 128:65 Util.scala 13:25]
  wire [15:0] _GEN_191 = _T_16 ? classmeta_reg_desc_state_field_type_13_sub_class_id : 16'h0; // @[Control.scala 126:39 Control.scala 128:65 Util.scala 13:25]
  wire [4:0] _GEN_192 = _T_16 ? classmeta_reg_desc_state_field_type_13_field_type : 5'h0; // @[Control.scala 126:39 Control.scala 128:65 Util.scala 13:25]
  wire  _GEN_193 = _T_16 & classmeta_reg_desc_state_field_type_13_is_repeated; // @[Control.scala 126:39 Control.scala 128:65 Util.scala 13:25]
  wire  _GEN_194 = _T_16 & classmeta_reg_desc_state_field_type_14_is_host; // @[Control.scala 126:39 Control.scala 128:65 Util.scala 13:25]
  wire [15:0] _GEN_195 = _T_16 ? classmeta_reg_desc_state_field_type_14_sub_class_id : 16'h0; // @[Control.scala 126:39 Control.scala 128:65 Util.scala 13:25]
  wire [4:0] _GEN_196 = _T_16 ? classmeta_reg_desc_state_field_type_14_field_type : 5'h0; // @[Control.scala 126:39 Control.scala 128:65 Util.scala 13:25]
  wire  _GEN_197 = _T_16 & classmeta_reg_desc_state_field_type_14_is_repeated; // @[Control.scala 126:39 Control.scala 128:65 Util.scala 13:25]
  wire  _GEN_198 = _T_16 & classmeta_reg_desc_state_field_type_15_is_host; // @[Control.scala 126:39 Control.scala 128:65 Util.scala 13:25]
  wire [15:0] _GEN_199 = _T_16 ? classmeta_reg_desc_state_field_type_15_sub_class_id : 16'h0; // @[Control.scala 126:39 Control.scala 128:65 Util.scala 13:25]
  wire [4:0] _GEN_200 = _T_16 ? classmeta_reg_desc_state_field_type_15_field_type : 5'h0; // @[Control.scala 126:39 Control.scala 128:65 Util.scala 13:25]
  wire  _GEN_201 = _T_16 & classmeta_reg_desc_state_field_type_15_is_repeated; // @[Control.scala 126:39 Control.scala 128:65 Util.scala 13:25]
  wire  _GEN_202 = _T_16 & classmeta_reg_desc_state_field_type_16_is_host; // @[Control.scala 126:39 Control.scala 128:65 Util.scala 13:25]
  wire [15:0] _GEN_203 = _T_16 ? classmeta_reg_desc_state_field_type_16_sub_class_id : 16'h0; // @[Control.scala 126:39 Control.scala 128:65 Util.scala 13:25]
  wire [4:0] _GEN_204 = _T_16 ? classmeta_reg_desc_state_field_type_16_field_type : 5'h0; // @[Control.scala 126:39 Control.scala 128:65 Util.scala 13:25]
  wire  _GEN_205 = _T_16 & classmeta_reg_desc_state_field_type_16_is_repeated; // @[Control.scala 126:39 Control.scala 128:65 Util.scala 13:25]
  wire  _GEN_206 = _T_16 & classmeta_reg_desc_state_field_type_17_is_host; // @[Control.scala 126:39 Control.scala 128:65 Util.scala 13:25]
  wire [15:0] _GEN_207 = _T_16 ? classmeta_reg_desc_state_field_type_17_sub_class_id : 16'h0; // @[Control.scala 126:39 Control.scala 128:65 Util.scala 13:25]
  wire [4:0] _GEN_208 = _T_16 ? classmeta_reg_desc_state_field_type_17_field_type : 5'h0; // @[Control.scala 126:39 Control.scala 128:65 Util.scala 13:25]
  wire  _GEN_209 = _T_16 & classmeta_reg_desc_state_field_type_17_is_repeated; // @[Control.scala 126:39 Control.scala 128:65 Util.scala 13:25]
  wire  _GEN_210 = _T_16 & classmeta_reg_desc_state_field_type_18_is_host; // @[Control.scala 126:39 Control.scala 128:65 Util.scala 13:25]
  wire [15:0] _GEN_211 = _T_16 ? classmeta_reg_desc_state_field_type_18_sub_class_id : 16'h0; // @[Control.scala 126:39 Control.scala 128:65 Util.scala 13:25]
  wire [4:0] _GEN_212 = _T_16 ? classmeta_reg_desc_state_field_type_18_field_type : 5'h0; // @[Control.scala 126:39 Control.scala 128:65 Util.scala 13:25]
  wire  _GEN_213 = _T_16 & classmeta_reg_desc_state_field_type_18_is_repeated; // @[Control.scala 126:39 Control.scala 128:65 Util.scala 13:25]
  wire  _GEN_214 = _T_16 & classmeta_reg_desc_state_field_type_19_is_host; // @[Control.scala 126:39 Control.scala 128:65 Util.scala 13:25]
  wire [15:0] _GEN_215 = _T_16 ? classmeta_reg_desc_state_field_type_19_sub_class_id : 16'h0; // @[Control.scala 126:39 Control.scala 128:65 Util.scala 13:25]
  wire [4:0] _GEN_216 = _T_16 ? classmeta_reg_desc_state_field_type_19_field_type : 5'h0; // @[Control.scala 126:39 Control.scala 128:65 Util.scala 13:25]
  wire  _GEN_217 = _T_16 & classmeta_reg_desc_state_field_type_19_is_repeated; // @[Control.scala 126:39 Control.scala 128:65 Util.scala 13:25]
  wire  _GEN_218 = _T_16 & classmeta_reg_desc_state_field_type_20_is_host; // @[Control.scala 126:39 Control.scala 128:65 Util.scala 13:25]
  wire [15:0] _GEN_219 = _T_16 ? classmeta_reg_desc_state_field_type_20_sub_class_id : 16'h0; // @[Control.scala 126:39 Control.scala 128:65 Util.scala 13:25]
  wire [4:0] _GEN_220 = _T_16 ? classmeta_reg_desc_state_field_type_20_field_type : 5'h0; // @[Control.scala 126:39 Control.scala 128:65 Util.scala 13:25]
  wire  _GEN_221 = _T_16 & classmeta_reg_desc_state_field_type_20_is_repeated; // @[Control.scala 126:39 Control.scala 128:65 Util.scala 13:25]
  wire  _GEN_222 = _T_16 & classmeta_reg_desc_state_field_type_21_is_host; // @[Control.scala 126:39 Control.scala 128:65 Util.scala 13:25]
  wire [15:0] _GEN_223 = _T_16 ? classmeta_reg_desc_state_field_type_21_sub_class_id : 16'h0; // @[Control.scala 126:39 Control.scala 128:65 Util.scala 13:25]
  wire [4:0] _GEN_224 = _T_16 ? classmeta_reg_desc_state_field_type_21_field_type : 5'h0; // @[Control.scala 126:39 Control.scala 128:65 Util.scala 13:25]
  wire  _GEN_225 = _T_16 & classmeta_reg_desc_state_field_type_21_is_repeated; // @[Control.scala 126:39 Control.scala 128:65 Util.scala 13:25]
  wire  _GEN_226 = _T_16 & classmeta_reg_desc_state_field_type_22_is_host; // @[Control.scala 126:39 Control.scala 128:65 Util.scala 13:25]
  wire [15:0] _GEN_227 = _T_16 ? classmeta_reg_desc_state_field_type_22_sub_class_id : 16'h0; // @[Control.scala 126:39 Control.scala 128:65 Util.scala 13:25]
  wire [4:0] _GEN_228 = _T_16 ? classmeta_reg_desc_state_field_type_22_field_type : 5'h0; // @[Control.scala 126:39 Control.scala 128:65 Util.scala 13:25]
  wire  _GEN_229 = _T_16 & classmeta_reg_desc_state_field_type_22_is_repeated; // @[Control.scala 126:39 Control.scala 128:65 Util.scala 13:25]
  wire  _GEN_230 = _T_16 & classmeta_reg_desc_state_field_type_23_is_host; // @[Control.scala 126:39 Control.scala 128:65 Util.scala 13:25]
  wire [15:0] _GEN_231 = _T_16 ? classmeta_reg_desc_state_field_type_23_sub_class_id : 16'h0; // @[Control.scala 126:39 Control.scala 128:65 Util.scala 13:25]
  wire [4:0] _GEN_232 = _T_16 ? classmeta_reg_desc_state_field_type_23_field_type : 5'h0; // @[Control.scala 126:39 Control.scala 128:65 Util.scala 13:25]
  wire  _GEN_233 = _T_16 & classmeta_reg_desc_state_field_type_23_is_repeated; // @[Control.scala 126:39 Control.scala 128:65 Util.scala 13:25]
  wire  _GEN_234 = _T_16 & classmeta_reg_desc_state_field_type_24_is_host; // @[Control.scala 126:39 Control.scala 128:65 Util.scala 13:25]
  wire [15:0] _GEN_235 = _T_16 ? classmeta_reg_desc_state_field_type_24_sub_class_id : 16'h0; // @[Control.scala 126:39 Control.scala 128:65 Util.scala 13:25]
  wire [4:0] _GEN_236 = _T_16 ? classmeta_reg_desc_state_field_type_24_field_type : 5'h0; // @[Control.scala 126:39 Control.scala 128:65 Util.scala 13:25]
  wire  _GEN_237 = _T_16 & classmeta_reg_desc_state_field_type_24_is_repeated; // @[Control.scala 126:39 Control.scala 128:65 Util.scala 13:25]
  wire  _GEN_238 = _T_16 & classmeta_reg_desc_state_field_type_25_is_host; // @[Control.scala 126:39 Control.scala 128:65 Util.scala 13:25]
  wire [15:0] _GEN_239 = _T_16 ? classmeta_reg_desc_state_field_type_25_sub_class_id : 16'h0; // @[Control.scala 126:39 Control.scala 128:65 Util.scala 13:25]
  wire [4:0] _GEN_240 = _T_16 ? classmeta_reg_desc_state_field_type_25_field_type : 5'h0; // @[Control.scala 126:39 Control.scala 128:65 Util.scala 13:25]
  wire  _GEN_241 = _T_16 & classmeta_reg_desc_state_field_type_25_is_repeated; // @[Control.scala 126:39 Control.scala 128:65 Util.scala 13:25]
  wire  _GEN_242 = _T_16 & classmeta_reg_desc_state_field_type_26_is_host; // @[Control.scala 126:39 Control.scala 128:65 Util.scala 13:25]
  wire [15:0] _GEN_243 = _T_16 ? classmeta_reg_desc_state_field_type_26_sub_class_id : 16'h0; // @[Control.scala 126:39 Control.scala 128:65 Util.scala 13:25]
  wire [4:0] _GEN_244 = _T_16 ? classmeta_reg_desc_state_field_type_26_field_type : 5'h0; // @[Control.scala 126:39 Control.scala 128:65 Util.scala 13:25]
  wire  _GEN_245 = _T_16 & classmeta_reg_desc_state_field_type_26_is_repeated; // @[Control.scala 126:39 Control.scala 128:65 Util.scala 13:25]
  wire  _GEN_246 = _T_16 & classmeta_reg_desc_state_field_type_27_is_host; // @[Control.scala 126:39 Control.scala 128:65 Util.scala 13:25]
  wire [15:0] _GEN_247 = _T_16 ? classmeta_reg_desc_state_field_type_27_sub_class_id : 16'h0; // @[Control.scala 126:39 Control.scala 128:65 Util.scala 13:25]
  wire [4:0] _GEN_248 = _T_16 ? classmeta_reg_desc_state_field_type_27_field_type : 5'h0; // @[Control.scala 126:39 Control.scala 128:65 Util.scala 13:25]
  wire  _GEN_249 = _T_16 & classmeta_reg_desc_state_field_type_27_is_repeated; // @[Control.scala 126:39 Control.scala 128:65 Util.scala 13:25]
  wire  _GEN_250 = _T_16 & classmeta_reg_desc_state_field_type_28_is_host; // @[Control.scala 126:39 Control.scala 128:65 Util.scala 13:25]
  wire [15:0] _GEN_251 = _T_16 ? classmeta_reg_desc_state_field_type_28_sub_class_id : 16'h0; // @[Control.scala 126:39 Control.scala 128:65 Util.scala 13:25]
  wire [4:0] _GEN_252 = _T_16 ? classmeta_reg_desc_state_field_type_28_field_type : 5'h0; // @[Control.scala 126:39 Control.scala 128:65 Util.scala 13:25]
  wire  _GEN_253 = _T_16 & classmeta_reg_desc_state_field_type_28_is_repeated; // @[Control.scala 126:39 Control.scala 128:65 Util.scala 13:25]
  wire  _GEN_254 = _T_16 & classmeta_reg_desc_state_field_type_29_is_host; // @[Control.scala 126:39 Control.scala 128:65 Util.scala 13:25]
  wire [15:0] _GEN_255 = _T_16 ? classmeta_reg_desc_state_field_type_29_sub_class_id : 16'h0; // @[Control.scala 126:39 Control.scala 128:65 Util.scala 13:25]
  wire [4:0] _GEN_256 = _T_16 ? classmeta_reg_desc_state_field_type_29_field_type : 5'h0; // @[Control.scala 126:39 Control.scala 128:65 Util.scala 13:25]
  wire  _GEN_257 = _T_16 & classmeta_reg_desc_state_field_type_29_is_repeated; // @[Control.scala 126:39 Control.scala 128:65 Util.scala 13:25]
  wire  _GEN_258 = _T_16 & io_axi_w_bits_data[0]; // @[Control.scala 126:39 Control.scala 131:84 Util.scala 13:25]
  wire [15:0] _GEN_259 = _T_16 ? io_axi_w_bits_data[31:16] : 16'h0; // @[Control.scala 126:39 Control.scala 134:84 Util.scala 13:25]
  wire [4:0] _GEN_260 = _T_16 ? io_axi_w_bits_data[6:2] : 5'h0; // @[Control.scala 126:39 Control.scala 133:84 Util.scala 13:25]
  wire  _GEN_261 = _T_16 & io_axi_w_bits_data[1]; // @[Control.scala 126:39 Control.scala 132:84 Util.scala 13:25]
  wire  _GEN_262 = _T_16 & io_axi_w_bits_data[32]; // @[Control.scala 126:39 Control.scala 131:84 Util.scala 13:25]
  wire [15:0] _GEN_263 = _T_16 ? io_axi_w_bits_data[63:48] : 16'h0; // @[Control.scala 126:39 Control.scala 134:84 Util.scala 13:25]
  wire [4:0] _GEN_264 = _T_16 ? io_axi_w_bits_data[38:34] : 5'h0; // @[Control.scala 126:39 Control.scala 133:84 Util.scala 13:25]
  wire  _GEN_265 = _T_16 & io_axi_w_bits_data[33]; // @[Control.scala 126:39 Control.scala 132:84 Util.scala 13:25]
  wire  _GEN_266 = _T_16 & io_axi_w_bits_data[64]; // @[Control.scala 126:39 Control.scala 131:84 Util.scala 13:25]
  wire [15:0] _GEN_267 = _T_16 ? io_axi_w_bits_data[95:80] : 16'h0; // @[Control.scala 126:39 Control.scala 134:84 Util.scala 13:25]
  wire [4:0] _GEN_268 = _T_16 ? io_axi_w_bits_data[70:66] : 5'h0; // @[Control.scala 126:39 Control.scala 133:84 Util.scala 13:25]
  wire  _GEN_269 = _T_16 & io_axi_w_bits_data[65]; // @[Control.scala 126:39 Control.scala 132:84 Util.scala 13:25]
  wire [7:0] _GEN_270 = _T_16 ? classmeta_reg_desc_state_max_field_num : 8'h0; // @[Control.scala 126:39 Control.scala 128:65 Util.scala 13:25]
  wire [15:0] _GEN_271 = _T_16 ? classmeta_reg_desc_state_class_length : 16'h0; // @[Control.scala 126:39 Control.scala 128:65 Util.scala 13:25]
  wire [9:0] _GEN_272 = _T_16 ? classmeta_reg_class_id : 10'h0; // @[Control.scala 126:39 Control.scala 128:65 Util.scala 13:25]
  wire  _GEN_273 = _T_16 ? 1'h0 : classmeta_reg_desc_state_field_type_0_is_host; // @[Control.scala 126:39 Control.scala 129:89 Control.scala 57:36]
  wire [15:0] _GEN_274 = _T_16 ? 16'h0 : classmeta_reg_desc_state_field_type_0_sub_class_id; // @[Control.scala 126:39 Control.scala 129:89 Control.scala 57:36]
  wire [4:0] _GEN_275 = _T_16 ? 5'h0 : classmeta_reg_desc_state_field_type_0_field_type; // @[Control.scala 126:39 Control.scala 129:89 Control.scala 57:36]
  wire  _GEN_276 = _T_16 ? 1'h0 : classmeta_reg_desc_state_field_type_0_is_repeated; // @[Control.scala 126:39 Control.scala 129:89 Control.scala 57:36]
  wire  _GEN_277 = _T_16 ? 1'h0 : classmeta_reg_desc_state_field_type_1_is_host; // @[Control.scala 126:39 Control.scala 129:89 Control.scala 57:36]
  wire [15:0] _GEN_278 = _T_16 ? 16'h0 : classmeta_reg_desc_state_field_type_1_sub_class_id; // @[Control.scala 126:39 Control.scala 129:89 Control.scala 57:36]
  wire [4:0] _GEN_279 = _T_16 ? 5'h0 : classmeta_reg_desc_state_field_type_1_field_type; // @[Control.scala 126:39 Control.scala 129:89 Control.scala 57:36]
  wire  _GEN_280 = _T_16 ? 1'h0 : classmeta_reg_desc_state_field_type_1_is_repeated; // @[Control.scala 126:39 Control.scala 129:89 Control.scala 57:36]
  wire  _GEN_281 = _T_16 ? 1'h0 : classmeta_reg_desc_state_field_type_2_is_host; // @[Control.scala 126:39 Control.scala 129:89 Control.scala 57:36]
  wire [15:0] _GEN_282 = _T_16 ? 16'h0 : classmeta_reg_desc_state_field_type_2_sub_class_id; // @[Control.scala 126:39 Control.scala 129:89 Control.scala 57:36]
  wire [4:0] _GEN_283 = _T_16 ? 5'h0 : classmeta_reg_desc_state_field_type_2_field_type; // @[Control.scala 126:39 Control.scala 129:89 Control.scala 57:36]
  wire  _GEN_284 = _T_16 ? 1'h0 : classmeta_reg_desc_state_field_type_2_is_repeated; // @[Control.scala 126:39 Control.scala 129:89 Control.scala 57:36]
  wire  _GEN_285 = _T_16 ? 1'h0 : classmeta_reg_desc_state_field_type_3_is_host; // @[Control.scala 126:39 Control.scala 129:89 Control.scala 57:36]
  wire [15:0] _GEN_286 = _T_16 ? 16'h0 : classmeta_reg_desc_state_field_type_3_sub_class_id; // @[Control.scala 126:39 Control.scala 129:89 Control.scala 57:36]
  wire [4:0] _GEN_287 = _T_16 ? 5'h0 : classmeta_reg_desc_state_field_type_3_field_type; // @[Control.scala 126:39 Control.scala 129:89 Control.scala 57:36]
  wire  _GEN_288 = _T_16 ? 1'h0 : classmeta_reg_desc_state_field_type_3_is_repeated; // @[Control.scala 126:39 Control.scala 129:89 Control.scala 57:36]
  wire  _GEN_289 = _T_16 ? 1'h0 : classmeta_reg_desc_state_field_type_4_is_host; // @[Control.scala 126:39 Control.scala 129:89 Control.scala 57:36]
  wire [15:0] _GEN_290 = _T_16 ? 16'h0 : classmeta_reg_desc_state_field_type_4_sub_class_id; // @[Control.scala 126:39 Control.scala 129:89 Control.scala 57:36]
  wire [4:0] _GEN_291 = _T_16 ? 5'h0 : classmeta_reg_desc_state_field_type_4_field_type; // @[Control.scala 126:39 Control.scala 129:89 Control.scala 57:36]
  wire  _GEN_292 = _T_16 ? 1'h0 : classmeta_reg_desc_state_field_type_4_is_repeated; // @[Control.scala 126:39 Control.scala 129:89 Control.scala 57:36]
  wire  _GEN_293 = _T_16 ? 1'h0 : classmeta_reg_desc_state_field_type_5_is_host; // @[Control.scala 126:39 Control.scala 129:89 Control.scala 57:36]
  wire [15:0] _GEN_294 = _T_16 ? 16'h0 : classmeta_reg_desc_state_field_type_5_sub_class_id; // @[Control.scala 126:39 Control.scala 129:89 Control.scala 57:36]
  wire [4:0] _GEN_295 = _T_16 ? 5'h0 : classmeta_reg_desc_state_field_type_5_field_type; // @[Control.scala 126:39 Control.scala 129:89 Control.scala 57:36]
  wire  _GEN_296 = _T_16 ? 1'h0 : classmeta_reg_desc_state_field_type_5_is_repeated; // @[Control.scala 126:39 Control.scala 129:89 Control.scala 57:36]
  wire  _GEN_297 = _T_16 ? 1'h0 : classmeta_reg_desc_state_field_type_6_is_host; // @[Control.scala 126:39 Control.scala 129:89 Control.scala 57:36]
  wire [15:0] _GEN_298 = _T_16 ? 16'h0 : classmeta_reg_desc_state_field_type_6_sub_class_id; // @[Control.scala 126:39 Control.scala 129:89 Control.scala 57:36]
  wire [4:0] _GEN_299 = _T_16 ? 5'h0 : classmeta_reg_desc_state_field_type_6_field_type; // @[Control.scala 126:39 Control.scala 129:89 Control.scala 57:36]
  wire  _GEN_300 = _T_16 ? 1'h0 : classmeta_reg_desc_state_field_type_6_is_repeated; // @[Control.scala 126:39 Control.scala 129:89 Control.scala 57:36]
  wire  _GEN_301 = _T_16 ? 1'h0 : classmeta_reg_desc_state_field_type_7_is_host; // @[Control.scala 126:39 Control.scala 129:89 Control.scala 57:36]
  wire [15:0] _GEN_302 = _T_16 ? 16'h0 : classmeta_reg_desc_state_field_type_7_sub_class_id; // @[Control.scala 126:39 Control.scala 129:89 Control.scala 57:36]
  wire [4:0] _GEN_303 = _T_16 ? 5'h0 : classmeta_reg_desc_state_field_type_7_field_type; // @[Control.scala 126:39 Control.scala 129:89 Control.scala 57:36]
  wire  _GEN_304 = _T_16 ? 1'h0 : classmeta_reg_desc_state_field_type_7_is_repeated; // @[Control.scala 126:39 Control.scala 129:89 Control.scala 57:36]
  wire  _GEN_305 = _T_16 ? 1'h0 : classmeta_reg_desc_state_field_type_8_is_host; // @[Control.scala 126:39 Control.scala 129:89 Control.scala 57:36]
  wire [15:0] _GEN_306 = _T_16 ? 16'h0 : classmeta_reg_desc_state_field_type_8_sub_class_id; // @[Control.scala 126:39 Control.scala 129:89 Control.scala 57:36]
  wire [4:0] _GEN_307 = _T_16 ? 5'h0 : classmeta_reg_desc_state_field_type_8_field_type; // @[Control.scala 126:39 Control.scala 129:89 Control.scala 57:36]
  wire  _GEN_308 = _T_16 ? 1'h0 : classmeta_reg_desc_state_field_type_8_is_repeated; // @[Control.scala 126:39 Control.scala 129:89 Control.scala 57:36]
  wire  _GEN_309 = _T_16 ? 1'h0 : classmeta_reg_desc_state_field_type_9_is_host; // @[Control.scala 126:39 Control.scala 129:89 Control.scala 57:36]
  wire [15:0] _GEN_310 = _T_16 ? 16'h0 : classmeta_reg_desc_state_field_type_9_sub_class_id; // @[Control.scala 126:39 Control.scala 129:89 Control.scala 57:36]
  wire [4:0] _GEN_311 = _T_16 ? 5'h0 : classmeta_reg_desc_state_field_type_9_field_type; // @[Control.scala 126:39 Control.scala 129:89 Control.scala 57:36]
  wire  _GEN_312 = _T_16 ? 1'h0 : classmeta_reg_desc_state_field_type_9_is_repeated; // @[Control.scala 126:39 Control.scala 129:89 Control.scala 57:36]
  wire  _GEN_313 = _T_16 ? 1'h0 : classmeta_reg_desc_state_field_type_10_is_host; // @[Control.scala 126:39 Control.scala 129:89 Control.scala 57:36]
  wire [15:0] _GEN_314 = _T_16 ? 16'h0 : classmeta_reg_desc_state_field_type_10_sub_class_id; // @[Control.scala 126:39 Control.scala 129:89 Control.scala 57:36]
  wire [4:0] _GEN_315 = _T_16 ? 5'h0 : classmeta_reg_desc_state_field_type_10_field_type; // @[Control.scala 126:39 Control.scala 129:89 Control.scala 57:36]
  wire  _GEN_316 = _T_16 ? 1'h0 : classmeta_reg_desc_state_field_type_10_is_repeated; // @[Control.scala 126:39 Control.scala 129:89 Control.scala 57:36]
  wire  _GEN_317 = _T_16 ? 1'h0 : classmeta_reg_desc_state_field_type_11_is_host; // @[Control.scala 126:39 Control.scala 129:89 Control.scala 57:36]
  wire [15:0] _GEN_318 = _T_16 ? 16'h0 : classmeta_reg_desc_state_field_type_11_sub_class_id; // @[Control.scala 126:39 Control.scala 129:89 Control.scala 57:36]
  wire [4:0] _GEN_319 = _T_16 ? 5'h0 : classmeta_reg_desc_state_field_type_11_field_type; // @[Control.scala 126:39 Control.scala 129:89 Control.scala 57:36]
  wire  _GEN_320 = _T_16 ? 1'h0 : classmeta_reg_desc_state_field_type_11_is_repeated; // @[Control.scala 126:39 Control.scala 129:89 Control.scala 57:36]
  wire  _GEN_321 = _T_16 ? 1'h0 : classmeta_reg_desc_state_field_type_12_is_host; // @[Control.scala 126:39 Control.scala 129:89 Control.scala 57:36]
  wire [15:0] _GEN_322 = _T_16 ? 16'h0 : classmeta_reg_desc_state_field_type_12_sub_class_id; // @[Control.scala 126:39 Control.scala 129:89 Control.scala 57:36]
  wire [4:0] _GEN_323 = _T_16 ? 5'h0 : classmeta_reg_desc_state_field_type_12_field_type; // @[Control.scala 126:39 Control.scala 129:89 Control.scala 57:36]
  wire  _GEN_324 = _T_16 ? 1'h0 : classmeta_reg_desc_state_field_type_12_is_repeated; // @[Control.scala 126:39 Control.scala 129:89 Control.scala 57:36]
  wire  _GEN_325 = _T_16 ? 1'h0 : classmeta_reg_desc_state_field_type_13_is_host; // @[Control.scala 126:39 Control.scala 129:89 Control.scala 57:36]
  wire [15:0] _GEN_326 = _T_16 ? 16'h0 : classmeta_reg_desc_state_field_type_13_sub_class_id; // @[Control.scala 126:39 Control.scala 129:89 Control.scala 57:36]
  wire [4:0] _GEN_327 = _T_16 ? 5'h0 : classmeta_reg_desc_state_field_type_13_field_type; // @[Control.scala 126:39 Control.scala 129:89 Control.scala 57:36]
  wire  _GEN_328 = _T_16 ? 1'h0 : classmeta_reg_desc_state_field_type_13_is_repeated; // @[Control.scala 126:39 Control.scala 129:89 Control.scala 57:36]
  wire  _GEN_329 = _T_16 ? 1'h0 : classmeta_reg_desc_state_field_type_14_is_host; // @[Control.scala 126:39 Control.scala 129:89 Control.scala 57:36]
  wire [15:0] _GEN_330 = _T_16 ? 16'h0 : classmeta_reg_desc_state_field_type_14_sub_class_id; // @[Control.scala 126:39 Control.scala 129:89 Control.scala 57:36]
  wire [4:0] _GEN_331 = _T_16 ? 5'h0 : classmeta_reg_desc_state_field_type_14_field_type; // @[Control.scala 126:39 Control.scala 129:89 Control.scala 57:36]
  wire  _GEN_332 = _T_16 ? 1'h0 : classmeta_reg_desc_state_field_type_14_is_repeated; // @[Control.scala 126:39 Control.scala 129:89 Control.scala 57:36]
  wire  _GEN_333 = _T_16 ? 1'h0 : classmeta_reg_desc_state_field_type_15_is_host; // @[Control.scala 126:39 Control.scala 129:89 Control.scala 57:36]
  wire [15:0] _GEN_334 = _T_16 ? 16'h0 : classmeta_reg_desc_state_field_type_15_sub_class_id; // @[Control.scala 126:39 Control.scala 129:89 Control.scala 57:36]
  wire [4:0] _GEN_335 = _T_16 ? 5'h0 : classmeta_reg_desc_state_field_type_15_field_type; // @[Control.scala 126:39 Control.scala 129:89 Control.scala 57:36]
  wire  _GEN_336 = _T_16 ? 1'h0 : classmeta_reg_desc_state_field_type_15_is_repeated; // @[Control.scala 126:39 Control.scala 129:89 Control.scala 57:36]
  wire  _GEN_337 = _T_16 ? 1'h0 : classmeta_reg_desc_state_field_type_16_is_host; // @[Control.scala 126:39 Control.scala 129:89 Control.scala 57:36]
  wire [15:0] _GEN_338 = _T_16 ? 16'h0 : classmeta_reg_desc_state_field_type_16_sub_class_id; // @[Control.scala 126:39 Control.scala 129:89 Control.scala 57:36]
  wire [4:0] _GEN_339 = _T_16 ? 5'h0 : classmeta_reg_desc_state_field_type_16_field_type; // @[Control.scala 126:39 Control.scala 129:89 Control.scala 57:36]
  wire  _GEN_340 = _T_16 ? 1'h0 : classmeta_reg_desc_state_field_type_16_is_repeated; // @[Control.scala 126:39 Control.scala 129:89 Control.scala 57:36]
  wire  _GEN_341 = _T_16 ? 1'h0 : classmeta_reg_desc_state_field_type_17_is_host; // @[Control.scala 126:39 Control.scala 129:89 Control.scala 57:36]
  wire [15:0] _GEN_342 = _T_16 ? 16'h0 : classmeta_reg_desc_state_field_type_17_sub_class_id; // @[Control.scala 126:39 Control.scala 129:89 Control.scala 57:36]
  wire [4:0] _GEN_343 = _T_16 ? 5'h0 : classmeta_reg_desc_state_field_type_17_field_type; // @[Control.scala 126:39 Control.scala 129:89 Control.scala 57:36]
  wire  _GEN_344 = _T_16 ? 1'h0 : classmeta_reg_desc_state_field_type_17_is_repeated; // @[Control.scala 126:39 Control.scala 129:89 Control.scala 57:36]
  wire  _GEN_345 = _T_16 ? 1'h0 : classmeta_reg_desc_state_field_type_18_is_host; // @[Control.scala 126:39 Control.scala 129:89 Control.scala 57:36]
  wire [15:0] _GEN_346 = _T_16 ? 16'h0 : classmeta_reg_desc_state_field_type_18_sub_class_id; // @[Control.scala 126:39 Control.scala 129:89 Control.scala 57:36]
  wire [4:0] _GEN_347 = _T_16 ? 5'h0 : classmeta_reg_desc_state_field_type_18_field_type; // @[Control.scala 126:39 Control.scala 129:89 Control.scala 57:36]
  wire  _GEN_348 = _T_16 ? 1'h0 : classmeta_reg_desc_state_field_type_18_is_repeated; // @[Control.scala 126:39 Control.scala 129:89 Control.scala 57:36]
  wire  _GEN_349 = _T_16 ? 1'h0 : classmeta_reg_desc_state_field_type_19_is_host; // @[Control.scala 126:39 Control.scala 129:89 Control.scala 57:36]
  wire [15:0] _GEN_350 = _T_16 ? 16'h0 : classmeta_reg_desc_state_field_type_19_sub_class_id; // @[Control.scala 126:39 Control.scala 129:89 Control.scala 57:36]
  wire [4:0] _GEN_351 = _T_16 ? 5'h0 : classmeta_reg_desc_state_field_type_19_field_type; // @[Control.scala 126:39 Control.scala 129:89 Control.scala 57:36]
  wire  _GEN_352 = _T_16 ? 1'h0 : classmeta_reg_desc_state_field_type_19_is_repeated; // @[Control.scala 126:39 Control.scala 129:89 Control.scala 57:36]
  wire  _GEN_353 = _T_16 ? 1'h0 : classmeta_reg_desc_state_field_type_20_is_host; // @[Control.scala 126:39 Control.scala 129:89 Control.scala 57:36]
  wire [15:0] _GEN_354 = _T_16 ? 16'h0 : classmeta_reg_desc_state_field_type_20_sub_class_id; // @[Control.scala 126:39 Control.scala 129:89 Control.scala 57:36]
  wire [4:0] _GEN_355 = _T_16 ? 5'h0 : classmeta_reg_desc_state_field_type_20_field_type; // @[Control.scala 126:39 Control.scala 129:89 Control.scala 57:36]
  wire  _GEN_356 = _T_16 ? 1'h0 : classmeta_reg_desc_state_field_type_20_is_repeated; // @[Control.scala 126:39 Control.scala 129:89 Control.scala 57:36]
  wire  _GEN_357 = _T_16 ? 1'h0 : classmeta_reg_desc_state_field_type_21_is_host; // @[Control.scala 126:39 Control.scala 129:89 Control.scala 57:36]
  wire [15:0] _GEN_358 = _T_16 ? 16'h0 : classmeta_reg_desc_state_field_type_21_sub_class_id; // @[Control.scala 126:39 Control.scala 129:89 Control.scala 57:36]
  wire [4:0] _GEN_359 = _T_16 ? 5'h0 : classmeta_reg_desc_state_field_type_21_field_type; // @[Control.scala 126:39 Control.scala 129:89 Control.scala 57:36]
  wire  _GEN_360 = _T_16 ? 1'h0 : classmeta_reg_desc_state_field_type_21_is_repeated; // @[Control.scala 126:39 Control.scala 129:89 Control.scala 57:36]
  wire  _GEN_361 = _T_16 ? 1'h0 : classmeta_reg_desc_state_field_type_22_is_host; // @[Control.scala 126:39 Control.scala 129:89 Control.scala 57:36]
  wire [15:0] _GEN_362 = _T_16 ? 16'h0 : classmeta_reg_desc_state_field_type_22_sub_class_id; // @[Control.scala 126:39 Control.scala 129:89 Control.scala 57:36]
  wire [4:0] _GEN_363 = _T_16 ? 5'h0 : classmeta_reg_desc_state_field_type_22_field_type; // @[Control.scala 126:39 Control.scala 129:89 Control.scala 57:36]
  wire  _GEN_364 = _T_16 ? 1'h0 : classmeta_reg_desc_state_field_type_22_is_repeated; // @[Control.scala 126:39 Control.scala 129:89 Control.scala 57:36]
  wire  _GEN_365 = _T_16 ? 1'h0 : classmeta_reg_desc_state_field_type_23_is_host; // @[Control.scala 126:39 Control.scala 129:89 Control.scala 57:36]
  wire [15:0] _GEN_366 = _T_16 ? 16'h0 : classmeta_reg_desc_state_field_type_23_sub_class_id; // @[Control.scala 126:39 Control.scala 129:89 Control.scala 57:36]
  wire [4:0] _GEN_367 = _T_16 ? 5'h0 : classmeta_reg_desc_state_field_type_23_field_type; // @[Control.scala 126:39 Control.scala 129:89 Control.scala 57:36]
  wire  _GEN_368 = _T_16 ? 1'h0 : classmeta_reg_desc_state_field_type_23_is_repeated; // @[Control.scala 126:39 Control.scala 129:89 Control.scala 57:36]
  wire  _GEN_369 = _T_16 ? 1'h0 : classmeta_reg_desc_state_field_type_24_is_host; // @[Control.scala 126:39 Control.scala 129:89 Control.scala 57:36]
  wire [15:0] _GEN_370 = _T_16 ? 16'h0 : classmeta_reg_desc_state_field_type_24_sub_class_id; // @[Control.scala 126:39 Control.scala 129:89 Control.scala 57:36]
  wire [4:0] _GEN_371 = _T_16 ? 5'h0 : classmeta_reg_desc_state_field_type_24_field_type; // @[Control.scala 126:39 Control.scala 129:89 Control.scala 57:36]
  wire  _GEN_372 = _T_16 ? 1'h0 : classmeta_reg_desc_state_field_type_24_is_repeated; // @[Control.scala 126:39 Control.scala 129:89 Control.scala 57:36]
  wire  _GEN_373 = _T_16 ? 1'h0 : classmeta_reg_desc_state_field_type_25_is_host; // @[Control.scala 126:39 Control.scala 129:89 Control.scala 57:36]
  wire [15:0] _GEN_374 = _T_16 ? 16'h0 : classmeta_reg_desc_state_field_type_25_sub_class_id; // @[Control.scala 126:39 Control.scala 129:89 Control.scala 57:36]
  wire [4:0] _GEN_375 = _T_16 ? 5'h0 : classmeta_reg_desc_state_field_type_25_field_type; // @[Control.scala 126:39 Control.scala 129:89 Control.scala 57:36]
  wire  _GEN_376 = _T_16 ? 1'h0 : classmeta_reg_desc_state_field_type_25_is_repeated; // @[Control.scala 126:39 Control.scala 129:89 Control.scala 57:36]
  wire  _GEN_377 = _T_16 ? 1'h0 : classmeta_reg_desc_state_field_type_26_is_host; // @[Control.scala 126:39 Control.scala 129:89 Control.scala 57:36]
  wire [15:0] _GEN_378 = _T_16 ? 16'h0 : classmeta_reg_desc_state_field_type_26_sub_class_id; // @[Control.scala 126:39 Control.scala 129:89 Control.scala 57:36]
  wire [4:0] _GEN_379 = _T_16 ? 5'h0 : classmeta_reg_desc_state_field_type_26_field_type; // @[Control.scala 126:39 Control.scala 129:89 Control.scala 57:36]
  wire  _GEN_380 = _T_16 ? 1'h0 : classmeta_reg_desc_state_field_type_26_is_repeated; // @[Control.scala 126:39 Control.scala 129:89 Control.scala 57:36]
  wire  _GEN_381 = _T_16 ? 1'h0 : classmeta_reg_desc_state_field_type_27_is_host; // @[Control.scala 126:39 Control.scala 129:89 Control.scala 57:36]
  wire [15:0] _GEN_382 = _T_16 ? 16'h0 : classmeta_reg_desc_state_field_type_27_sub_class_id; // @[Control.scala 126:39 Control.scala 129:89 Control.scala 57:36]
  wire [4:0] _GEN_383 = _T_16 ? 5'h0 : classmeta_reg_desc_state_field_type_27_field_type; // @[Control.scala 126:39 Control.scala 129:89 Control.scala 57:36]
  wire  _GEN_384 = _T_16 ? 1'h0 : classmeta_reg_desc_state_field_type_27_is_repeated; // @[Control.scala 126:39 Control.scala 129:89 Control.scala 57:36]
  wire  _GEN_385 = _T_16 ? 1'h0 : classmeta_reg_desc_state_field_type_28_is_host; // @[Control.scala 126:39 Control.scala 129:89 Control.scala 57:36]
  wire [15:0] _GEN_386 = _T_16 ? 16'h0 : classmeta_reg_desc_state_field_type_28_sub_class_id; // @[Control.scala 126:39 Control.scala 129:89 Control.scala 57:36]
  wire [4:0] _GEN_387 = _T_16 ? 5'h0 : classmeta_reg_desc_state_field_type_28_field_type; // @[Control.scala 126:39 Control.scala 129:89 Control.scala 57:36]
  wire  _GEN_388 = _T_16 ? 1'h0 : classmeta_reg_desc_state_field_type_28_is_repeated; // @[Control.scala 126:39 Control.scala 129:89 Control.scala 57:36]
  wire  _GEN_389 = _T_16 ? 1'h0 : classmeta_reg_desc_state_field_type_29_is_host; // @[Control.scala 126:39 Control.scala 129:89 Control.scala 57:36]
  wire [15:0] _GEN_390 = _T_16 ? 16'h0 : classmeta_reg_desc_state_field_type_29_sub_class_id; // @[Control.scala 126:39 Control.scala 129:89 Control.scala 57:36]
  wire [4:0] _GEN_391 = _T_16 ? 5'h0 : classmeta_reg_desc_state_field_type_29_field_type; // @[Control.scala 126:39 Control.scala 129:89 Control.scala 57:36]
  wire  _GEN_392 = _T_16 ? 1'h0 : classmeta_reg_desc_state_field_type_29_is_repeated; // @[Control.scala 126:39 Control.scala 129:89 Control.scala 57:36]
  wire [7:0] _GEN_405 = _T_16 ? 8'h0 : classmeta_reg_desc_state_max_field_num; // @[Control.scala 126:39 Control.scala 129:89 Control.scala 57:36]
  wire [15:0] _GEN_406 = _T_16 ? 16'h0 : classmeta_reg_desc_state_class_length; // @[Control.scala 126:39 Control.scala 129:89 Control.scala 57:36]
  wire [9:0] _GEN_407 = _T_16 ? 10'h0 : classmeta_reg_class_id; // @[Control.scala 126:39 Control.scala 129:89 Control.scala 57:36]
  wire  _T_23 = 3'h6 == s_wr; // @[Conditional.scala 37:30]
  wire [10:0] _GEN_410 = _T_16 ? io_axi_w_bits_data[10:0] : 11'h0; // @[Control.scala 140:39 Control.scala 142:53 Util.scala 13:25]
  wire [63:0] _GEN_411 = _T_16 ? io_axi_w_bits_data[127:64] : 64'h0; // @[Control.scala 140:39 Control.scala 143:53 Util.scala 13:25]
  wire  _T_25 = 3'h7 == s_wr; // @[Conditional.scala 37:30]
  wire  _T_27 = 3'h1 == s_wr; // @[Conditional.scala 37:30]
  wire [2:0] _GEN_426 = _T_27 ? _GEN_11 : s_wr; // @[Conditional.scala 39:67 Control.scala 43:27]
  wire [2:0] _GEN_434 = _T_25 ? _GEN_11 : _GEN_426; // @[Conditional.scala 39:67]
  wire [10:0] _GEN_436 = _T_23 ? _GEN_410 : 11'h0; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [63:0] _GEN_437 = _T_23 ? _GEN_411 : 64'h0; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [2:0] _GEN_442 = _T_23 ? _GEN_11 : _GEN_434; // @[Conditional.scala 39:67]
  wire [15:0] _GEN_452 = _T_21 ? _GEN_139 : 16'h0; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [4:0] _GEN_453 = _T_21 ? _GEN_140 : 5'h0; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [15:0] _GEN_456 = _T_21 ? _GEN_143 : 16'h0; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [4:0] _GEN_457 = _T_21 ? _GEN_144 : 5'h0; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [15:0] _GEN_460 = _T_21 ? _GEN_147 : 16'h0; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [4:0] _GEN_461 = _T_21 ? _GEN_148 : 5'h0; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [15:0] _GEN_464 = _T_21 ? _GEN_151 : 16'h0; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [4:0] _GEN_465 = _T_21 ? _GEN_152 : 5'h0; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [15:0] _GEN_468 = _T_21 ? _GEN_155 : 16'h0; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [4:0] _GEN_469 = _T_21 ? _GEN_156 : 5'h0; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [15:0] _GEN_472 = _T_21 ? _GEN_159 : 16'h0; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [4:0] _GEN_473 = _T_21 ? _GEN_160 : 5'h0; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [15:0] _GEN_476 = _T_21 ? _GEN_163 : 16'h0; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [4:0] _GEN_477 = _T_21 ? _GEN_164 : 5'h0; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [15:0] _GEN_480 = _T_21 ? _GEN_167 : 16'h0; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [4:0] _GEN_481 = _T_21 ? _GEN_168 : 5'h0; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [15:0] _GEN_484 = _T_21 ? _GEN_171 : 16'h0; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [4:0] _GEN_485 = _T_21 ? _GEN_172 : 5'h0; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [15:0] _GEN_488 = _T_21 ? _GEN_175 : 16'h0; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [4:0] _GEN_489 = _T_21 ? _GEN_176 : 5'h0; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [15:0] _GEN_492 = _T_21 ? _GEN_179 : 16'h0; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [4:0] _GEN_493 = _T_21 ? _GEN_180 : 5'h0; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [15:0] _GEN_496 = _T_21 ? _GEN_183 : 16'h0; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [4:0] _GEN_497 = _T_21 ? _GEN_184 : 5'h0; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [15:0] _GEN_500 = _T_21 ? _GEN_187 : 16'h0; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [4:0] _GEN_501 = _T_21 ? _GEN_188 : 5'h0; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [15:0] _GEN_504 = _T_21 ? _GEN_191 : 16'h0; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [4:0] _GEN_505 = _T_21 ? _GEN_192 : 5'h0; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [15:0] _GEN_508 = _T_21 ? _GEN_195 : 16'h0; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [4:0] _GEN_509 = _T_21 ? _GEN_196 : 5'h0; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [15:0] _GEN_512 = _T_21 ? _GEN_199 : 16'h0; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [4:0] _GEN_513 = _T_21 ? _GEN_200 : 5'h0; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [15:0] _GEN_516 = _T_21 ? _GEN_203 : 16'h0; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [4:0] _GEN_517 = _T_21 ? _GEN_204 : 5'h0; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [15:0] _GEN_520 = _T_21 ? _GEN_207 : 16'h0; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [4:0] _GEN_521 = _T_21 ? _GEN_208 : 5'h0; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [15:0] _GEN_524 = _T_21 ? _GEN_211 : 16'h0; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [4:0] _GEN_525 = _T_21 ? _GEN_212 : 5'h0; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [15:0] _GEN_528 = _T_21 ? _GEN_215 : 16'h0; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [4:0] _GEN_529 = _T_21 ? _GEN_216 : 5'h0; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [15:0] _GEN_532 = _T_21 ? _GEN_219 : 16'h0; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [4:0] _GEN_533 = _T_21 ? _GEN_220 : 5'h0; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [15:0] _GEN_536 = _T_21 ? _GEN_223 : 16'h0; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [4:0] _GEN_537 = _T_21 ? _GEN_224 : 5'h0; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [15:0] _GEN_540 = _T_21 ? _GEN_227 : 16'h0; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [4:0] _GEN_541 = _T_21 ? _GEN_228 : 5'h0; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [15:0] _GEN_544 = _T_21 ? _GEN_231 : 16'h0; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [4:0] _GEN_545 = _T_21 ? _GEN_232 : 5'h0; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [15:0] _GEN_548 = _T_21 ? _GEN_235 : 16'h0; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [4:0] _GEN_549 = _T_21 ? _GEN_236 : 5'h0; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [15:0] _GEN_552 = _T_21 ? _GEN_239 : 16'h0; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [4:0] _GEN_553 = _T_21 ? _GEN_240 : 5'h0; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [15:0] _GEN_556 = _T_21 ? _GEN_243 : 16'h0; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [4:0] _GEN_557 = _T_21 ? _GEN_244 : 5'h0; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [15:0] _GEN_560 = _T_21 ? _GEN_247 : 16'h0; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [4:0] _GEN_561 = _T_21 ? _GEN_248 : 5'h0; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [15:0] _GEN_564 = _T_21 ? _GEN_251 : 16'h0; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [4:0] _GEN_565 = _T_21 ? _GEN_252 : 5'h0; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [15:0] _GEN_568 = _T_21 ? _GEN_255 : 16'h0; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [4:0] _GEN_569 = _T_21 ? _GEN_256 : 5'h0; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [15:0] _GEN_572 = _T_21 ? _GEN_259 : 16'h0; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [4:0] _GEN_573 = _T_21 ? _GEN_260 : 5'h0; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [15:0] _GEN_576 = _T_21 ? _GEN_263 : 16'h0; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [4:0] _GEN_577 = _T_21 ? _GEN_264 : 5'h0; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [15:0] _GEN_580 = _T_21 ? _GEN_267 : 16'h0; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [4:0] _GEN_581 = _T_21 ? _GEN_268 : 5'h0; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [7:0] _GEN_583 = _T_21 ? _GEN_270 : 8'h0; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [15:0] _GEN_584 = _T_21 ? _GEN_271 : 16'h0; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [9:0] _GEN_585 = _T_21 ? _GEN_272 : 10'h0; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire  _GEN_586 = _T_21 ? _GEN_273 : classmeta_reg_desc_state_field_type_0_is_host; // @[Conditional.scala 39:67 Control.scala 57:36]
  wire [15:0] _GEN_587 = _T_21 ? _GEN_274 : classmeta_reg_desc_state_field_type_0_sub_class_id; // @[Conditional.scala 39:67 Control.scala 57:36]
  wire [4:0] _GEN_588 = _T_21 ? _GEN_275 : classmeta_reg_desc_state_field_type_0_field_type; // @[Conditional.scala 39:67 Control.scala 57:36]
  wire  _GEN_589 = _T_21 ? _GEN_276 : classmeta_reg_desc_state_field_type_0_is_repeated; // @[Conditional.scala 39:67 Control.scala 57:36]
  wire  _GEN_590 = _T_21 ? _GEN_277 : classmeta_reg_desc_state_field_type_1_is_host; // @[Conditional.scala 39:67 Control.scala 57:36]
  wire [15:0] _GEN_591 = _T_21 ? _GEN_278 : classmeta_reg_desc_state_field_type_1_sub_class_id; // @[Conditional.scala 39:67 Control.scala 57:36]
  wire [4:0] _GEN_592 = _T_21 ? _GEN_279 : classmeta_reg_desc_state_field_type_1_field_type; // @[Conditional.scala 39:67 Control.scala 57:36]
  wire  _GEN_593 = _T_21 ? _GEN_280 : classmeta_reg_desc_state_field_type_1_is_repeated; // @[Conditional.scala 39:67 Control.scala 57:36]
  wire  _GEN_594 = _T_21 ? _GEN_281 : classmeta_reg_desc_state_field_type_2_is_host; // @[Conditional.scala 39:67 Control.scala 57:36]
  wire [15:0] _GEN_595 = _T_21 ? _GEN_282 : classmeta_reg_desc_state_field_type_2_sub_class_id; // @[Conditional.scala 39:67 Control.scala 57:36]
  wire [4:0] _GEN_596 = _T_21 ? _GEN_283 : classmeta_reg_desc_state_field_type_2_field_type; // @[Conditional.scala 39:67 Control.scala 57:36]
  wire  _GEN_597 = _T_21 ? _GEN_284 : classmeta_reg_desc_state_field_type_2_is_repeated; // @[Conditional.scala 39:67 Control.scala 57:36]
  wire  _GEN_598 = _T_21 ? _GEN_285 : classmeta_reg_desc_state_field_type_3_is_host; // @[Conditional.scala 39:67 Control.scala 57:36]
  wire [15:0] _GEN_599 = _T_21 ? _GEN_286 : classmeta_reg_desc_state_field_type_3_sub_class_id; // @[Conditional.scala 39:67 Control.scala 57:36]
  wire [4:0] _GEN_600 = _T_21 ? _GEN_287 : classmeta_reg_desc_state_field_type_3_field_type; // @[Conditional.scala 39:67 Control.scala 57:36]
  wire  _GEN_601 = _T_21 ? _GEN_288 : classmeta_reg_desc_state_field_type_3_is_repeated; // @[Conditional.scala 39:67 Control.scala 57:36]
  wire  _GEN_602 = _T_21 ? _GEN_289 : classmeta_reg_desc_state_field_type_4_is_host; // @[Conditional.scala 39:67 Control.scala 57:36]
  wire [15:0] _GEN_603 = _T_21 ? _GEN_290 : classmeta_reg_desc_state_field_type_4_sub_class_id; // @[Conditional.scala 39:67 Control.scala 57:36]
  wire [4:0] _GEN_604 = _T_21 ? _GEN_291 : classmeta_reg_desc_state_field_type_4_field_type; // @[Conditional.scala 39:67 Control.scala 57:36]
  wire  _GEN_605 = _T_21 ? _GEN_292 : classmeta_reg_desc_state_field_type_4_is_repeated; // @[Conditional.scala 39:67 Control.scala 57:36]
  wire  _GEN_606 = _T_21 ? _GEN_293 : classmeta_reg_desc_state_field_type_5_is_host; // @[Conditional.scala 39:67 Control.scala 57:36]
  wire [15:0] _GEN_607 = _T_21 ? _GEN_294 : classmeta_reg_desc_state_field_type_5_sub_class_id; // @[Conditional.scala 39:67 Control.scala 57:36]
  wire [4:0] _GEN_608 = _T_21 ? _GEN_295 : classmeta_reg_desc_state_field_type_5_field_type; // @[Conditional.scala 39:67 Control.scala 57:36]
  wire  _GEN_609 = _T_21 ? _GEN_296 : classmeta_reg_desc_state_field_type_5_is_repeated; // @[Conditional.scala 39:67 Control.scala 57:36]
  wire  _GEN_610 = _T_21 ? _GEN_297 : classmeta_reg_desc_state_field_type_6_is_host; // @[Conditional.scala 39:67 Control.scala 57:36]
  wire [15:0] _GEN_611 = _T_21 ? _GEN_298 : classmeta_reg_desc_state_field_type_6_sub_class_id; // @[Conditional.scala 39:67 Control.scala 57:36]
  wire [4:0] _GEN_612 = _T_21 ? _GEN_299 : classmeta_reg_desc_state_field_type_6_field_type; // @[Conditional.scala 39:67 Control.scala 57:36]
  wire  _GEN_613 = _T_21 ? _GEN_300 : classmeta_reg_desc_state_field_type_6_is_repeated; // @[Conditional.scala 39:67 Control.scala 57:36]
  wire  _GEN_614 = _T_21 ? _GEN_301 : classmeta_reg_desc_state_field_type_7_is_host; // @[Conditional.scala 39:67 Control.scala 57:36]
  wire [15:0] _GEN_615 = _T_21 ? _GEN_302 : classmeta_reg_desc_state_field_type_7_sub_class_id; // @[Conditional.scala 39:67 Control.scala 57:36]
  wire [4:0] _GEN_616 = _T_21 ? _GEN_303 : classmeta_reg_desc_state_field_type_7_field_type; // @[Conditional.scala 39:67 Control.scala 57:36]
  wire  _GEN_617 = _T_21 ? _GEN_304 : classmeta_reg_desc_state_field_type_7_is_repeated; // @[Conditional.scala 39:67 Control.scala 57:36]
  wire  _GEN_618 = _T_21 ? _GEN_305 : classmeta_reg_desc_state_field_type_8_is_host; // @[Conditional.scala 39:67 Control.scala 57:36]
  wire [15:0] _GEN_619 = _T_21 ? _GEN_306 : classmeta_reg_desc_state_field_type_8_sub_class_id; // @[Conditional.scala 39:67 Control.scala 57:36]
  wire [4:0] _GEN_620 = _T_21 ? _GEN_307 : classmeta_reg_desc_state_field_type_8_field_type; // @[Conditional.scala 39:67 Control.scala 57:36]
  wire  _GEN_621 = _T_21 ? _GEN_308 : classmeta_reg_desc_state_field_type_8_is_repeated; // @[Conditional.scala 39:67 Control.scala 57:36]
  wire  _GEN_622 = _T_21 ? _GEN_309 : classmeta_reg_desc_state_field_type_9_is_host; // @[Conditional.scala 39:67 Control.scala 57:36]
  wire [15:0] _GEN_623 = _T_21 ? _GEN_310 : classmeta_reg_desc_state_field_type_9_sub_class_id; // @[Conditional.scala 39:67 Control.scala 57:36]
  wire [4:0] _GEN_624 = _T_21 ? _GEN_311 : classmeta_reg_desc_state_field_type_9_field_type; // @[Conditional.scala 39:67 Control.scala 57:36]
  wire  _GEN_625 = _T_21 ? _GEN_312 : classmeta_reg_desc_state_field_type_9_is_repeated; // @[Conditional.scala 39:67 Control.scala 57:36]
  wire  _GEN_626 = _T_21 ? _GEN_313 : classmeta_reg_desc_state_field_type_10_is_host; // @[Conditional.scala 39:67 Control.scala 57:36]
  wire [15:0] _GEN_627 = _T_21 ? _GEN_314 : classmeta_reg_desc_state_field_type_10_sub_class_id; // @[Conditional.scala 39:67 Control.scala 57:36]
  wire [4:0] _GEN_628 = _T_21 ? _GEN_315 : classmeta_reg_desc_state_field_type_10_field_type; // @[Conditional.scala 39:67 Control.scala 57:36]
  wire  _GEN_629 = _T_21 ? _GEN_316 : classmeta_reg_desc_state_field_type_10_is_repeated; // @[Conditional.scala 39:67 Control.scala 57:36]
  wire  _GEN_630 = _T_21 ? _GEN_317 : classmeta_reg_desc_state_field_type_11_is_host; // @[Conditional.scala 39:67 Control.scala 57:36]
  wire [15:0] _GEN_631 = _T_21 ? _GEN_318 : classmeta_reg_desc_state_field_type_11_sub_class_id; // @[Conditional.scala 39:67 Control.scala 57:36]
  wire [4:0] _GEN_632 = _T_21 ? _GEN_319 : classmeta_reg_desc_state_field_type_11_field_type; // @[Conditional.scala 39:67 Control.scala 57:36]
  wire  _GEN_633 = _T_21 ? _GEN_320 : classmeta_reg_desc_state_field_type_11_is_repeated; // @[Conditional.scala 39:67 Control.scala 57:36]
  wire  _GEN_634 = _T_21 ? _GEN_321 : classmeta_reg_desc_state_field_type_12_is_host; // @[Conditional.scala 39:67 Control.scala 57:36]
  wire [15:0] _GEN_635 = _T_21 ? _GEN_322 : classmeta_reg_desc_state_field_type_12_sub_class_id; // @[Conditional.scala 39:67 Control.scala 57:36]
  wire [4:0] _GEN_636 = _T_21 ? _GEN_323 : classmeta_reg_desc_state_field_type_12_field_type; // @[Conditional.scala 39:67 Control.scala 57:36]
  wire  _GEN_637 = _T_21 ? _GEN_324 : classmeta_reg_desc_state_field_type_12_is_repeated; // @[Conditional.scala 39:67 Control.scala 57:36]
  wire  _GEN_638 = _T_21 ? _GEN_325 : classmeta_reg_desc_state_field_type_13_is_host; // @[Conditional.scala 39:67 Control.scala 57:36]
  wire [15:0] _GEN_639 = _T_21 ? _GEN_326 : classmeta_reg_desc_state_field_type_13_sub_class_id; // @[Conditional.scala 39:67 Control.scala 57:36]
  wire [4:0] _GEN_640 = _T_21 ? _GEN_327 : classmeta_reg_desc_state_field_type_13_field_type; // @[Conditional.scala 39:67 Control.scala 57:36]
  wire  _GEN_641 = _T_21 ? _GEN_328 : classmeta_reg_desc_state_field_type_13_is_repeated; // @[Conditional.scala 39:67 Control.scala 57:36]
  wire  _GEN_642 = _T_21 ? _GEN_329 : classmeta_reg_desc_state_field_type_14_is_host; // @[Conditional.scala 39:67 Control.scala 57:36]
  wire [15:0] _GEN_643 = _T_21 ? _GEN_330 : classmeta_reg_desc_state_field_type_14_sub_class_id; // @[Conditional.scala 39:67 Control.scala 57:36]
  wire [4:0] _GEN_644 = _T_21 ? _GEN_331 : classmeta_reg_desc_state_field_type_14_field_type; // @[Conditional.scala 39:67 Control.scala 57:36]
  wire  _GEN_645 = _T_21 ? _GEN_332 : classmeta_reg_desc_state_field_type_14_is_repeated; // @[Conditional.scala 39:67 Control.scala 57:36]
  wire  _GEN_646 = _T_21 ? _GEN_333 : classmeta_reg_desc_state_field_type_15_is_host; // @[Conditional.scala 39:67 Control.scala 57:36]
  wire [15:0] _GEN_647 = _T_21 ? _GEN_334 : classmeta_reg_desc_state_field_type_15_sub_class_id; // @[Conditional.scala 39:67 Control.scala 57:36]
  wire [4:0] _GEN_648 = _T_21 ? _GEN_335 : classmeta_reg_desc_state_field_type_15_field_type; // @[Conditional.scala 39:67 Control.scala 57:36]
  wire  _GEN_649 = _T_21 ? _GEN_336 : classmeta_reg_desc_state_field_type_15_is_repeated; // @[Conditional.scala 39:67 Control.scala 57:36]
  wire  _GEN_650 = _T_21 ? _GEN_337 : classmeta_reg_desc_state_field_type_16_is_host; // @[Conditional.scala 39:67 Control.scala 57:36]
  wire [15:0] _GEN_651 = _T_21 ? _GEN_338 : classmeta_reg_desc_state_field_type_16_sub_class_id; // @[Conditional.scala 39:67 Control.scala 57:36]
  wire [4:0] _GEN_652 = _T_21 ? _GEN_339 : classmeta_reg_desc_state_field_type_16_field_type; // @[Conditional.scala 39:67 Control.scala 57:36]
  wire  _GEN_653 = _T_21 ? _GEN_340 : classmeta_reg_desc_state_field_type_16_is_repeated; // @[Conditional.scala 39:67 Control.scala 57:36]
  wire  _GEN_654 = _T_21 ? _GEN_341 : classmeta_reg_desc_state_field_type_17_is_host; // @[Conditional.scala 39:67 Control.scala 57:36]
  wire [15:0] _GEN_655 = _T_21 ? _GEN_342 : classmeta_reg_desc_state_field_type_17_sub_class_id; // @[Conditional.scala 39:67 Control.scala 57:36]
  wire [4:0] _GEN_656 = _T_21 ? _GEN_343 : classmeta_reg_desc_state_field_type_17_field_type; // @[Conditional.scala 39:67 Control.scala 57:36]
  wire  _GEN_657 = _T_21 ? _GEN_344 : classmeta_reg_desc_state_field_type_17_is_repeated; // @[Conditional.scala 39:67 Control.scala 57:36]
  wire  _GEN_658 = _T_21 ? _GEN_345 : classmeta_reg_desc_state_field_type_18_is_host; // @[Conditional.scala 39:67 Control.scala 57:36]
  wire [15:0] _GEN_659 = _T_21 ? _GEN_346 : classmeta_reg_desc_state_field_type_18_sub_class_id; // @[Conditional.scala 39:67 Control.scala 57:36]
  wire [4:0] _GEN_660 = _T_21 ? _GEN_347 : classmeta_reg_desc_state_field_type_18_field_type; // @[Conditional.scala 39:67 Control.scala 57:36]
  wire  _GEN_661 = _T_21 ? _GEN_348 : classmeta_reg_desc_state_field_type_18_is_repeated; // @[Conditional.scala 39:67 Control.scala 57:36]
  wire  _GEN_662 = _T_21 ? _GEN_349 : classmeta_reg_desc_state_field_type_19_is_host; // @[Conditional.scala 39:67 Control.scala 57:36]
  wire [15:0] _GEN_663 = _T_21 ? _GEN_350 : classmeta_reg_desc_state_field_type_19_sub_class_id; // @[Conditional.scala 39:67 Control.scala 57:36]
  wire [4:0] _GEN_664 = _T_21 ? _GEN_351 : classmeta_reg_desc_state_field_type_19_field_type; // @[Conditional.scala 39:67 Control.scala 57:36]
  wire  _GEN_665 = _T_21 ? _GEN_352 : classmeta_reg_desc_state_field_type_19_is_repeated; // @[Conditional.scala 39:67 Control.scala 57:36]
  wire  _GEN_666 = _T_21 ? _GEN_353 : classmeta_reg_desc_state_field_type_20_is_host; // @[Conditional.scala 39:67 Control.scala 57:36]
  wire [15:0] _GEN_667 = _T_21 ? _GEN_354 : classmeta_reg_desc_state_field_type_20_sub_class_id; // @[Conditional.scala 39:67 Control.scala 57:36]
  wire [4:0] _GEN_668 = _T_21 ? _GEN_355 : classmeta_reg_desc_state_field_type_20_field_type; // @[Conditional.scala 39:67 Control.scala 57:36]
  wire  _GEN_669 = _T_21 ? _GEN_356 : classmeta_reg_desc_state_field_type_20_is_repeated; // @[Conditional.scala 39:67 Control.scala 57:36]
  wire  _GEN_670 = _T_21 ? _GEN_357 : classmeta_reg_desc_state_field_type_21_is_host; // @[Conditional.scala 39:67 Control.scala 57:36]
  wire [15:0] _GEN_671 = _T_21 ? _GEN_358 : classmeta_reg_desc_state_field_type_21_sub_class_id; // @[Conditional.scala 39:67 Control.scala 57:36]
  wire [4:0] _GEN_672 = _T_21 ? _GEN_359 : classmeta_reg_desc_state_field_type_21_field_type; // @[Conditional.scala 39:67 Control.scala 57:36]
  wire  _GEN_673 = _T_21 ? _GEN_360 : classmeta_reg_desc_state_field_type_21_is_repeated; // @[Conditional.scala 39:67 Control.scala 57:36]
  wire  _GEN_674 = _T_21 ? _GEN_361 : classmeta_reg_desc_state_field_type_22_is_host; // @[Conditional.scala 39:67 Control.scala 57:36]
  wire [15:0] _GEN_675 = _T_21 ? _GEN_362 : classmeta_reg_desc_state_field_type_22_sub_class_id; // @[Conditional.scala 39:67 Control.scala 57:36]
  wire [4:0] _GEN_676 = _T_21 ? _GEN_363 : classmeta_reg_desc_state_field_type_22_field_type; // @[Conditional.scala 39:67 Control.scala 57:36]
  wire  _GEN_677 = _T_21 ? _GEN_364 : classmeta_reg_desc_state_field_type_22_is_repeated; // @[Conditional.scala 39:67 Control.scala 57:36]
  wire  _GEN_678 = _T_21 ? _GEN_365 : classmeta_reg_desc_state_field_type_23_is_host; // @[Conditional.scala 39:67 Control.scala 57:36]
  wire [15:0] _GEN_679 = _T_21 ? _GEN_366 : classmeta_reg_desc_state_field_type_23_sub_class_id; // @[Conditional.scala 39:67 Control.scala 57:36]
  wire [4:0] _GEN_680 = _T_21 ? _GEN_367 : classmeta_reg_desc_state_field_type_23_field_type; // @[Conditional.scala 39:67 Control.scala 57:36]
  wire  _GEN_681 = _T_21 ? _GEN_368 : classmeta_reg_desc_state_field_type_23_is_repeated; // @[Conditional.scala 39:67 Control.scala 57:36]
  wire  _GEN_682 = _T_21 ? _GEN_369 : classmeta_reg_desc_state_field_type_24_is_host; // @[Conditional.scala 39:67 Control.scala 57:36]
  wire [15:0] _GEN_683 = _T_21 ? _GEN_370 : classmeta_reg_desc_state_field_type_24_sub_class_id; // @[Conditional.scala 39:67 Control.scala 57:36]
  wire [4:0] _GEN_684 = _T_21 ? _GEN_371 : classmeta_reg_desc_state_field_type_24_field_type; // @[Conditional.scala 39:67 Control.scala 57:36]
  wire  _GEN_685 = _T_21 ? _GEN_372 : classmeta_reg_desc_state_field_type_24_is_repeated; // @[Conditional.scala 39:67 Control.scala 57:36]
  wire  _GEN_686 = _T_21 ? _GEN_373 : classmeta_reg_desc_state_field_type_25_is_host; // @[Conditional.scala 39:67 Control.scala 57:36]
  wire [15:0] _GEN_687 = _T_21 ? _GEN_374 : classmeta_reg_desc_state_field_type_25_sub_class_id; // @[Conditional.scala 39:67 Control.scala 57:36]
  wire [4:0] _GEN_688 = _T_21 ? _GEN_375 : classmeta_reg_desc_state_field_type_25_field_type; // @[Conditional.scala 39:67 Control.scala 57:36]
  wire  _GEN_689 = _T_21 ? _GEN_376 : classmeta_reg_desc_state_field_type_25_is_repeated; // @[Conditional.scala 39:67 Control.scala 57:36]
  wire  _GEN_690 = _T_21 ? _GEN_377 : classmeta_reg_desc_state_field_type_26_is_host; // @[Conditional.scala 39:67 Control.scala 57:36]
  wire [15:0] _GEN_691 = _T_21 ? _GEN_378 : classmeta_reg_desc_state_field_type_26_sub_class_id; // @[Conditional.scala 39:67 Control.scala 57:36]
  wire [4:0] _GEN_692 = _T_21 ? _GEN_379 : classmeta_reg_desc_state_field_type_26_field_type; // @[Conditional.scala 39:67 Control.scala 57:36]
  wire  _GEN_693 = _T_21 ? _GEN_380 : classmeta_reg_desc_state_field_type_26_is_repeated; // @[Conditional.scala 39:67 Control.scala 57:36]
  wire  _GEN_694 = _T_21 ? _GEN_381 : classmeta_reg_desc_state_field_type_27_is_host; // @[Conditional.scala 39:67 Control.scala 57:36]
  wire [15:0] _GEN_695 = _T_21 ? _GEN_382 : classmeta_reg_desc_state_field_type_27_sub_class_id; // @[Conditional.scala 39:67 Control.scala 57:36]
  wire [4:0] _GEN_696 = _T_21 ? _GEN_383 : classmeta_reg_desc_state_field_type_27_field_type; // @[Conditional.scala 39:67 Control.scala 57:36]
  wire  _GEN_697 = _T_21 ? _GEN_384 : classmeta_reg_desc_state_field_type_27_is_repeated; // @[Conditional.scala 39:67 Control.scala 57:36]
  wire  _GEN_698 = _T_21 ? _GEN_385 : classmeta_reg_desc_state_field_type_28_is_host; // @[Conditional.scala 39:67 Control.scala 57:36]
  wire [15:0] _GEN_699 = _T_21 ? _GEN_386 : classmeta_reg_desc_state_field_type_28_sub_class_id; // @[Conditional.scala 39:67 Control.scala 57:36]
  wire [4:0] _GEN_700 = _T_21 ? _GEN_387 : classmeta_reg_desc_state_field_type_28_field_type; // @[Conditional.scala 39:67 Control.scala 57:36]
  wire  _GEN_701 = _T_21 ? _GEN_388 : classmeta_reg_desc_state_field_type_28_is_repeated; // @[Conditional.scala 39:67 Control.scala 57:36]
  wire  _GEN_702 = _T_21 ? _GEN_389 : classmeta_reg_desc_state_field_type_29_is_host; // @[Conditional.scala 39:67 Control.scala 57:36]
  wire [15:0] _GEN_703 = _T_21 ? _GEN_390 : classmeta_reg_desc_state_field_type_29_sub_class_id; // @[Conditional.scala 39:67 Control.scala 57:36]
  wire [4:0] _GEN_704 = _T_21 ? _GEN_391 : classmeta_reg_desc_state_field_type_29_field_type; // @[Conditional.scala 39:67 Control.scala 57:36]
  wire  _GEN_705 = _T_21 ? _GEN_392 : classmeta_reg_desc_state_field_type_29_is_repeated; // @[Conditional.scala 39:67 Control.scala 57:36]
  wire [7:0] _GEN_718 = _T_21 ? _GEN_405 : classmeta_reg_desc_state_max_field_num; // @[Conditional.scala 39:67 Control.scala 57:36]
  wire [15:0] _GEN_719 = _T_21 ? _GEN_406 : classmeta_reg_desc_state_class_length; // @[Conditional.scala 39:67 Control.scala 57:36]
  wire [9:0] _GEN_720 = _T_21 ? _GEN_407 : classmeta_reg_class_id; // @[Conditional.scala 39:67 Control.scala 57:36]
  wire [2:0] _GEN_721 = _T_21 ? _GEN_11 : _GEN_442; // @[Conditional.scala 39:67]
  wire  _GEN_722 = _T_21 ? 1'h0 : _T_23 & _T_16; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [10:0] _GEN_723 = _T_21 ? 11'h0 : _GEN_436; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [63:0] _GEN_724 = _T_21 ? 64'h0 : _GEN_437; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire  _GEN_736 = _T_19 ? _GEN_72 : _GEN_642; // @[Conditional.scala 39:67]
  wire  _GEN_737 = _T_19 ? _GEN_73 : _GEN_645; // @[Conditional.scala 39:67]
  wire [4:0] _GEN_738 = _T_19 ? _GEN_74 : _GEN_644; // @[Conditional.scala 39:67]
  wire [15:0] _GEN_739 = _T_19 ? _GEN_75 : _GEN_643; // @[Conditional.scala 39:67]
  wire  _GEN_740 = _T_19 ? _GEN_76 : _GEN_646; // @[Conditional.scala 39:67]
  wire  _GEN_741 = _T_19 ? _GEN_77 : _GEN_649; // @[Conditional.scala 39:67]
  wire [4:0] _GEN_742 = _T_19 ? _GEN_78 : _GEN_648; // @[Conditional.scala 39:67]
  wire [15:0] _GEN_743 = _T_19 ? _GEN_79 : _GEN_647; // @[Conditional.scala 39:67]
  wire  _GEN_744 = _T_19 ? _GEN_80 : _GEN_650; // @[Conditional.scala 39:67]
  wire  _GEN_745 = _T_19 ? _GEN_81 : _GEN_653; // @[Conditional.scala 39:67]
  wire [4:0] _GEN_746 = _T_19 ? _GEN_82 : _GEN_652; // @[Conditional.scala 39:67]
  wire [15:0] _GEN_747 = _T_19 ? _GEN_83 : _GEN_651; // @[Conditional.scala 39:67]
  wire  _GEN_748 = _T_19 ? _GEN_84 : _GEN_654; // @[Conditional.scala 39:67]
  wire  _GEN_749 = _T_19 ? _GEN_85 : _GEN_657; // @[Conditional.scala 39:67]
  wire [4:0] _GEN_750 = _T_19 ? _GEN_86 : _GEN_656; // @[Conditional.scala 39:67]
  wire [15:0] _GEN_751 = _T_19 ? _GEN_87 : _GEN_655; // @[Conditional.scala 39:67]
  wire  _GEN_752 = _T_19 ? _GEN_88 : _GEN_658; // @[Conditional.scala 39:67]
  wire  _GEN_753 = _T_19 ? _GEN_89 : _GEN_661; // @[Conditional.scala 39:67]
  wire [4:0] _GEN_754 = _T_19 ? _GEN_90 : _GEN_660; // @[Conditional.scala 39:67]
  wire [15:0] _GEN_755 = _T_19 ? _GEN_91 : _GEN_659; // @[Conditional.scala 39:67]
  wire  _GEN_756 = _T_19 ? _GEN_92 : _GEN_662; // @[Conditional.scala 39:67]
  wire  _GEN_757 = _T_19 ? _GEN_93 : _GEN_665; // @[Conditional.scala 39:67]
  wire [4:0] _GEN_758 = _T_19 ? _GEN_94 : _GEN_664; // @[Conditional.scala 39:67]
  wire [15:0] _GEN_759 = _T_19 ? _GEN_95 : _GEN_663; // @[Conditional.scala 39:67]
  wire  _GEN_760 = _T_19 ? _GEN_96 : _GEN_666; // @[Conditional.scala 39:67]
  wire  _GEN_761 = _T_19 ? _GEN_97 : _GEN_669; // @[Conditional.scala 39:67]
  wire [4:0] _GEN_762 = _T_19 ? _GEN_98 : _GEN_668; // @[Conditional.scala 39:67]
  wire [15:0] _GEN_763 = _T_19 ? _GEN_99 : _GEN_667; // @[Conditional.scala 39:67]
  wire  _GEN_764 = _T_19 ? _GEN_100 : _GEN_670; // @[Conditional.scala 39:67]
  wire  _GEN_765 = _T_19 ? _GEN_101 : _GEN_673; // @[Conditional.scala 39:67]
  wire [4:0] _GEN_766 = _T_19 ? _GEN_102 : _GEN_672; // @[Conditional.scala 39:67]
  wire [15:0] _GEN_767 = _T_19 ? _GEN_103 : _GEN_671; // @[Conditional.scala 39:67]
  wire  _GEN_768 = _T_19 ? _GEN_104 : _GEN_674; // @[Conditional.scala 39:67]
  wire  _GEN_769 = _T_19 ? _GEN_105 : _GEN_677; // @[Conditional.scala 39:67]
  wire [4:0] _GEN_770 = _T_19 ? _GEN_106 : _GEN_676; // @[Conditional.scala 39:67]
  wire [15:0] _GEN_771 = _T_19 ? _GEN_107 : _GEN_675; // @[Conditional.scala 39:67]
  wire  _GEN_772 = _T_19 ? _GEN_108 : _GEN_678; // @[Conditional.scala 39:67]
  wire  _GEN_773 = _T_19 ? _GEN_109 : _GEN_681; // @[Conditional.scala 39:67]
  wire [4:0] _GEN_774 = _T_19 ? _GEN_110 : _GEN_680; // @[Conditional.scala 39:67]
  wire [15:0] _GEN_775 = _T_19 ? _GEN_111 : _GEN_679; // @[Conditional.scala 39:67]
  wire  _GEN_776 = _T_19 ? _GEN_112 : _GEN_682; // @[Conditional.scala 39:67]
  wire  _GEN_777 = _T_19 ? _GEN_113 : _GEN_685; // @[Conditional.scala 39:67]
  wire [4:0] _GEN_778 = _T_19 ? _GEN_114 : _GEN_684; // @[Conditional.scala 39:67]
  wire [15:0] _GEN_779 = _T_19 ? _GEN_115 : _GEN_683; // @[Conditional.scala 39:67]
  wire  _GEN_780 = _T_19 ? _GEN_116 : _GEN_686; // @[Conditional.scala 39:67]
  wire  _GEN_781 = _T_19 ? _GEN_117 : _GEN_689; // @[Conditional.scala 39:67]
  wire [4:0] _GEN_782 = _T_19 ? _GEN_118 : _GEN_688; // @[Conditional.scala 39:67]
  wire [15:0] _GEN_783 = _T_19 ? _GEN_119 : _GEN_687; // @[Conditional.scala 39:67]
  wire  _GEN_784 = _T_19 ? _GEN_120 : _GEN_690; // @[Conditional.scala 39:67]
  wire  _GEN_785 = _T_19 ? _GEN_121 : _GEN_693; // @[Conditional.scala 39:67]
  wire [4:0] _GEN_786 = _T_19 ? _GEN_122 : _GEN_692; // @[Conditional.scala 39:67]
  wire [15:0] _GEN_787 = _T_19 ? _GEN_123 : _GEN_691; // @[Conditional.scala 39:67]
  wire  _GEN_788 = _T_19 ? _GEN_124 : _GEN_694; // @[Conditional.scala 39:67]
  wire  _GEN_789 = _T_19 ? _GEN_125 : _GEN_697; // @[Conditional.scala 39:67]
  wire [4:0] _GEN_790 = _T_19 ? _GEN_126 : _GEN_696; // @[Conditional.scala 39:67]
  wire [15:0] _GEN_791 = _T_19 ? _GEN_127 : _GEN_695; // @[Conditional.scala 39:67]
  wire  _GEN_792 = _T_19 ? _GEN_128 : _GEN_698; // @[Conditional.scala 39:67]
  wire  _GEN_793 = _T_19 ? _GEN_129 : _GEN_701; // @[Conditional.scala 39:67]
  wire [4:0] _GEN_794 = _T_19 ? _GEN_130 : _GEN_700; // @[Conditional.scala 39:67]
  wire [15:0] _GEN_795 = _T_19 ? _GEN_131 : _GEN_699; // @[Conditional.scala 39:67]
  wire  _GEN_796 = _T_19 ? _GEN_132 : _GEN_702; // @[Conditional.scala 39:67]
  wire  _GEN_797 = _T_19 ? _GEN_133 : _GEN_705; // @[Conditional.scala 39:67]
  wire [4:0] _GEN_798 = _T_19 ? _GEN_134 : _GEN_704; // @[Conditional.scala 39:67]
  wire [15:0] _GEN_799 = _T_19 ? _GEN_135 : _GEN_703; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_800 = _T_19 ? _GEN_11 : _GEN_721; // @[Conditional.scala 39:67]
  wire  _GEN_801 = _T_19 ? 1'h0 : _T_21 & _T_16; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire  _GEN_802 = _T_19 ? 1'h0 : _T_21 & _GEN_138; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [15:0] _GEN_803 = _T_19 ? 16'h0 : _GEN_452; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [4:0] _GEN_804 = _T_19 ? 5'h0 : _GEN_453; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire  _GEN_805 = _T_19 ? 1'h0 : _T_21 & _GEN_141; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire  _GEN_806 = _T_19 ? 1'h0 : _T_21 & _GEN_142; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [15:0] _GEN_807 = _T_19 ? 16'h0 : _GEN_456; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [4:0] _GEN_808 = _T_19 ? 5'h0 : _GEN_457; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire  _GEN_809 = _T_19 ? 1'h0 : _T_21 & _GEN_145; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire  _GEN_810 = _T_19 ? 1'h0 : _T_21 & _GEN_146; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [15:0] _GEN_811 = _T_19 ? 16'h0 : _GEN_460; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [4:0] _GEN_812 = _T_19 ? 5'h0 : _GEN_461; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire  _GEN_813 = _T_19 ? 1'h0 : _T_21 & _GEN_149; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire  _GEN_814 = _T_19 ? 1'h0 : _T_21 & _GEN_150; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [15:0] _GEN_815 = _T_19 ? 16'h0 : _GEN_464; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [4:0] _GEN_816 = _T_19 ? 5'h0 : _GEN_465; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire  _GEN_817 = _T_19 ? 1'h0 : _T_21 & _GEN_153; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire  _GEN_818 = _T_19 ? 1'h0 : _T_21 & _GEN_154; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [15:0] _GEN_819 = _T_19 ? 16'h0 : _GEN_468; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [4:0] _GEN_820 = _T_19 ? 5'h0 : _GEN_469; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire  _GEN_821 = _T_19 ? 1'h0 : _T_21 & _GEN_157; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire  _GEN_822 = _T_19 ? 1'h0 : _T_21 & _GEN_158; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [15:0] _GEN_823 = _T_19 ? 16'h0 : _GEN_472; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [4:0] _GEN_824 = _T_19 ? 5'h0 : _GEN_473; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire  _GEN_825 = _T_19 ? 1'h0 : _T_21 & _GEN_161; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire  _GEN_826 = _T_19 ? 1'h0 : _T_21 & _GEN_162; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [15:0] _GEN_827 = _T_19 ? 16'h0 : _GEN_476; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [4:0] _GEN_828 = _T_19 ? 5'h0 : _GEN_477; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire  _GEN_829 = _T_19 ? 1'h0 : _T_21 & _GEN_165; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire  _GEN_830 = _T_19 ? 1'h0 : _T_21 & _GEN_166; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [15:0] _GEN_831 = _T_19 ? 16'h0 : _GEN_480; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [4:0] _GEN_832 = _T_19 ? 5'h0 : _GEN_481; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire  _GEN_833 = _T_19 ? 1'h0 : _T_21 & _GEN_169; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire  _GEN_834 = _T_19 ? 1'h0 : _T_21 & _GEN_170; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [15:0] _GEN_835 = _T_19 ? 16'h0 : _GEN_484; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [4:0] _GEN_836 = _T_19 ? 5'h0 : _GEN_485; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire  _GEN_837 = _T_19 ? 1'h0 : _T_21 & _GEN_173; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire  _GEN_838 = _T_19 ? 1'h0 : _T_21 & _GEN_174; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [15:0] _GEN_839 = _T_19 ? 16'h0 : _GEN_488; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [4:0] _GEN_840 = _T_19 ? 5'h0 : _GEN_489; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire  _GEN_841 = _T_19 ? 1'h0 : _T_21 & _GEN_177; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire  _GEN_842 = _T_19 ? 1'h0 : _T_21 & _GEN_178; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [15:0] _GEN_843 = _T_19 ? 16'h0 : _GEN_492; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [4:0] _GEN_844 = _T_19 ? 5'h0 : _GEN_493; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire  _GEN_845 = _T_19 ? 1'h0 : _T_21 & _GEN_181; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire  _GEN_846 = _T_19 ? 1'h0 : _T_21 & _GEN_182; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [15:0] _GEN_847 = _T_19 ? 16'h0 : _GEN_496; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [4:0] _GEN_848 = _T_19 ? 5'h0 : _GEN_497; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire  _GEN_849 = _T_19 ? 1'h0 : _T_21 & _GEN_185; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire  _GEN_850 = _T_19 ? 1'h0 : _T_21 & _GEN_186; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [15:0] _GEN_851 = _T_19 ? 16'h0 : _GEN_500; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [4:0] _GEN_852 = _T_19 ? 5'h0 : _GEN_501; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire  _GEN_853 = _T_19 ? 1'h0 : _T_21 & _GEN_189; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire  _GEN_854 = _T_19 ? 1'h0 : _T_21 & _GEN_190; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [15:0] _GEN_855 = _T_19 ? 16'h0 : _GEN_504; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [4:0] _GEN_856 = _T_19 ? 5'h0 : _GEN_505; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire  _GEN_857 = _T_19 ? 1'h0 : _T_21 & _GEN_193; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire  _GEN_858 = _T_19 ? 1'h0 : _T_21 & _GEN_194; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [15:0] _GEN_859 = _T_19 ? 16'h0 : _GEN_508; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [4:0] _GEN_860 = _T_19 ? 5'h0 : _GEN_509; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire  _GEN_861 = _T_19 ? 1'h0 : _T_21 & _GEN_197; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire  _GEN_862 = _T_19 ? 1'h0 : _T_21 & _GEN_198; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [15:0] _GEN_863 = _T_19 ? 16'h0 : _GEN_512; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [4:0] _GEN_864 = _T_19 ? 5'h0 : _GEN_513; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire  _GEN_865 = _T_19 ? 1'h0 : _T_21 & _GEN_201; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire  _GEN_866 = _T_19 ? 1'h0 : _T_21 & _GEN_202; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [15:0] _GEN_867 = _T_19 ? 16'h0 : _GEN_516; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [4:0] _GEN_868 = _T_19 ? 5'h0 : _GEN_517; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire  _GEN_869 = _T_19 ? 1'h0 : _T_21 & _GEN_205; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire  _GEN_870 = _T_19 ? 1'h0 : _T_21 & _GEN_206; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [15:0] _GEN_871 = _T_19 ? 16'h0 : _GEN_520; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [4:0] _GEN_872 = _T_19 ? 5'h0 : _GEN_521; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire  _GEN_873 = _T_19 ? 1'h0 : _T_21 & _GEN_209; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire  _GEN_874 = _T_19 ? 1'h0 : _T_21 & _GEN_210; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [15:0] _GEN_875 = _T_19 ? 16'h0 : _GEN_524; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [4:0] _GEN_876 = _T_19 ? 5'h0 : _GEN_525; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire  _GEN_877 = _T_19 ? 1'h0 : _T_21 & _GEN_213; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire  _GEN_878 = _T_19 ? 1'h0 : _T_21 & _GEN_214; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [15:0] _GEN_879 = _T_19 ? 16'h0 : _GEN_528; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [4:0] _GEN_880 = _T_19 ? 5'h0 : _GEN_529; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire  _GEN_881 = _T_19 ? 1'h0 : _T_21 & _GEN_217; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire  _GEN_882 = _T_19 ? 1'h0 : _T_21 & _GEN_218; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [15:0] _GEN_883 = _T_19 ? 16'h0 : _GEN_532; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [4:0] _GEN_884 = _T_19 ? 5'h0 : _GEN_533; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire  _GEN_885 = _T_19 ? 1'h0 : _T_21 & _GEN_221; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire  _GEN_886 = _T_19 ? 1'h0 : _T_21 & _GEN_222; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [15:0] _GEN_887 = _T_19 ? 16'h0 : _GEN_536; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [4:0] _GEN_888 = _T_19 ? 5'h0 : _GEN_537; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire  _GEN_889 = _T_19 ? 1'h0 : _T_21 & _GEN_225; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire  _GEN_890 = _T_19 ? 1'h0 : _T_21 & _GEN_226; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [15:0] _GEN_891 = _T_19 ? 16'h0 : _GEN_540; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [4:0] _GEN_892 = _T_19 ? 5'h0 : _GEN_541; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire  _GEN_893 = _T_19 ? 1'h0 : _T_21 & _GEN_229; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire  _GEN_894 = _T_19 ? 1'h0 : _T_21 & _GEN_230; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [15:0] _GEN_895 = _T_19 ? 16'h0 : _GEN_544; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [4:0] _GEN_896 = _T_19 ? 5'h0 : _GEN_545; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire  _GEN_897 = _T_19 ? 1'h0 : _T_21 & _GEN_233; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire  _GEN_898 = _T_19 ? 1'h0 : _T_21 & _GEN_234; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [15:0] _GEN_899 = _T_19 ? 16'h0 : _GEN_548; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [4:0] _GEN_900 = _T_19 ? 5'h0 : _GEN_549; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire  _GEN_901 = _T_19 ? 1'h0 : _T_21 & _GEN_237; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire  _GEN_902 = _T_19 ? 1'h0 : _T_21 & _GEN_238; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [15:0] _GEN_903 = _T_19 ? 16'h0 : _GEN_552; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [4:0] _GEN_904 = _T_19 ? 5'h0 : _GEN_553; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire  _GEN_905 = _T_19 ? 1'h0 : _T_21 & _GEN_241; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire  _GEN_906 = _T_19 ? 1'h0 : _T_21 & _GEN_242; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [15:0] _GEN_907 = _T_19 ? 16'h0 : _GEN_556; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [4:0] _GEN_908 = _T_19 ? 5'h0 : _GEN_557; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire  _GEN_909 = _T_19 ? 1'h0 : _T_21 & _GEN_245; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire  _GEN_910 = _T_19 ? 1'h0 : _T_21 & _GEN_246; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [15:0] _GEN_911 = _T_19 ? 16'h0 : _GEN_560; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [4:0] _GEN_912 = _T_19 ? 5'h0 : _GEN_561; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire  _GEN_913 = _T_19 ? 1'h0 : _T_21 & _GEN_249; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire  _GEN_914 = _T_19 ? 1'h0 : _T_21 & _GEN_250; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [15:0] _GEN_915 = _T_19 ? 16'h0 : _GEN_564; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [4:0] _GEN_916 = _T_19 ? 5'h0 : _GEN_565; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire  _GEN_917 = _T_19 ? 1'h0 : _T_21 & _GEN_253; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire  _GEN_918 = _T_19 ? 1'h0 : _T_21 & _GEN_254; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [15:0] _GEN_919 = _T_19 ? 16'h0 : _GEN_568; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [4:0] _GEN_920 = _T_19 ? 5'h0 : _GEN_569; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire  _GEN_921 = _T_19 ? 1'h0 : _T_21 & _GEN_257; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire  _GEN_922 = _T_19 ? 1'h0 : _T_21 & _GEN_258; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [15:0] _GEN_923 = _T_19 ? 16'h0 : _GEN_572; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [4:0] _GEN_924 = _T_19 ? 5'h0 : _GEN_573; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire  _GEN_925 = _T_19 ? 1'h0 : _T_21 & _GEN_261; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire  _GEN_926 = _T_19 ? 1'h0 : _T_21 & _GEN_262; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [15:0] _GEN_927 = _T_19 ? 16'h0 : _GEN_576; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [4:0] _GEN_928 = _T_19 ? 5'h0 : _GEN_577; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire  _GEN_929 = _T_19 ? 1'h0 : _T_21 & _GEN_265; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire  _GEN_930 = _T_19 ? 1'h0 : _T_21 & _GEN_266; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [15:0] _GEN_931 = _T_19 ? 16'h0 : _GEN_580; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [4:0] _GEN_932 = _T_19 ? 5'h0 : _GEN_581; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire  _GEN_933 = _T_19 ? 1'h0 : _T_21 & _GEN_269; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [7:0] _GEN_934 = _T_19 ? 8'h0 : _GEN_583; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [15:0] _GEN_935 = _T_19 ? 16'h0 : _GEN_584; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [9:0] _GEN_936 = _T_19 ? 10'h0 : _GEN_585; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire  _GEN_937 = _T_19 ? classmeta_reg_desc_state_field_type_0_is_host : _GEN_586; // @[Conditional.scala 39:67 Control.scala 57:36]
  wire [15:0] _GEN_938 = _T_19 ? classmeta_reg_desc_state_field_type_0_sub_class_id : _GEN_587; // @[Conditional.scala 39:67 Control.scala 57:36]
  wire [4:0] _GEN_939 = _T_19 ? classmeta_reg_desc_state_field_type_0_field_type : _GEN_588; // @[Conditional.scala 39:67 Control.scala 57:36]
  wire  _GEN_940 = _T_19 ? classmeta_reg_desc_state_field_type_0_is_repeated : _GEN_589; // @[Conditional.scala 39:67 Control.scala 57:36]
  wire  _GEN_941 = _T_19 ? classmeta_reg_desc_state_field_type_1_is_host : _GEN_590; // @[Conditional.scala 39:67 Control.scala 57:36]
  wire [15:0] _GEN_942 = _T_19 ? classmeta_reg_desc_state_field_type_1_sub_class_id : _GEN_591; // @[Conditional.scala 39:67 Control.scala 57:36]
  wire [4:0] _GEN_943 = _T_19 ? classmeta_reg_desc_state_field_type_1_field_type : _GEN_592; // @[Conditional.scala 39:67 Control.scala 57:36]
  wire  _GEN_944 = _T_19 ? classmeta_reg_desc_state_field_type_1_is_repeated : _GEN_593; // @[Conditional.scala 39:67 Control.scala 57:36]
  wire  _GEN_945 = _T_19 ? classmeta_reg_desc_state_field_type_2_is_host : _GEN_594; // @[Conditional.scala 39:67 Control.scala 57:36]
  wire [15:0] _GEN_946 = _T_19 ? classmeta_reg_desc_state_field_type_2_sub_class_id : _GEN_595; // @[Conditional.scala 39:67 Control.scala 57:36]
  wire [4:0] _GEN_947 = _T_19 ? classmeta_reg_desc_state_field_type_2_field_type : _GEN_596; // @[Conditional.scala 39:67 Control.scala 57:36]
  wire  _GEN_948 = _T_19 ? classmeta_reg_desc_state_field_type_2_is_repeated : _GEN_597; // @[Conditional.scala 39:67 Control.scala 57:36]
  wire  _GEN_949 = _T_19 ? classmeta_reg_desc_state_field_type_3_is_host : _GEN_598; // @[Conditional.scala 39:67 Control.scala 57:36]
  wire [15:0] _GEN_950 = _T_19 ? classmeta_reg_desc_state_field_type_3_sub_class_id : _GEN_599; // @[Conditional.scala 39:67 Control.scala 57:36]
  wire [4:0] _GEN_951 = _T_19 ? classmeta_reg_desc_state_field_type_3_field_type : _GEN_600; // @[Conditional.scala 39:67 Control.scala 57:36]
  wire  _GEN_952 = _T_19 ? classmeta_reg_desc_state_field_type_3_is_repeated : _GEN_601; // @[Conditional.scala 39:67 Control.scala 57:36]
  wire  _GEN_953 = _T_19 ? classmeta_reg_desc_state_field_type_4_is_host : _GEN_602; // @[Conditional.scala 39:67 Control.scala 57:36]
  wire [15:0] _GEN_954 = _T_19 ? classmeta_reg_desc_state_field_type_4_sub_class_id : _GEN_603; // @[Conditional.scala 39:67 Control.scala 57:36]
  wire [4:0] _GEN_955 = _T_19 ? classmeta_reg_desc_state_field_type_4_field_type : _GEN_604; // @[Conditional.scala 39:67 Control.scala 57:36]
  wire  _GEN_956 = _T_19 ? classmeta_reg_desc_state_field_type_4_is_repeated : _GEN_605; // @[Conditional.scala 39:67 Control.scala 57:36]
  wire  _GEN_957 = _T_19 ? classmeta_reg_desc_state_field_type_5_is_host : _GEN_606; // @[Conditional.scala 39:67 Control.scala 57:36]
  wire [15:0] _GEN_958 = _T_19 ? classmeta_reg_desc_state_field_type_5_sub_class_id : _GEN_607; // @[Conditional.scala 39:67 Control.scala 57:36]
  wire [4:0] _GEN_959 = _T_19 ? classmeta_reg_desc_state_field_type_5_field_type : _GEN_608; // @[Conditional.scala 39:67 Control.scala 57:36]
  wire  _GEN_960 = _T_19 ? classmeta_reg_desc_state_field_type_5_is_repeated : _GEN_609; // @[Conditional.scala 39:67 Control.scala 57:36]
  wire  _GEN_961 = _T_19 ? classmeta_reg_desc_state_field_type_6_is_host : _GEN_610; // @[Conditional.scala 39:67 Control.scala 57:36]
  wire [15:0] _GEN_962 = _T_19 ? classmeta_reg_desc_state_field_type_6_sub_class_id : _GEN_611; // @[Conditional.scala 39:67 Control.scala 57:36]
  wire [4:0] _GEN_963 = _T_19 ? classmeta_reg_desc_state_field_type_6_field_type : _GEN_612; // @[Conditional.scala 39:67 Control.scala 57:36]
  wire  _GEN_964 = _T_19 ? classmeta_reg_desc_state_field_type_6_is_repeated : _GEN_613; // @[Conditional.scala 39:67 Control.scala 57:36]
  wire  _GEN_965 = _T_19 ? classmeta_reg_desc_state_field_type_7_is_host : _GEN_614; // @[Conditional.scala 39:67 Control.scala 57:36]
  wire [15:0] _GEN_966 = _T_19 ? classmeta_reg_desc_state_field_type_7_sub_class_id : _GEN_615; // @[Conditional.scala 39:67 Control.scala 57:36]
  wire [4:0] _GEN_967 = _T_19 ? classmeta_reg_desc_state_field_type_7_field_type : _GEN_616; // @[Conditional.scala 39:67 Control.scala 57:36]
  wire  _GEN_968 = _T_19 ? classmeta_reg_desc_state_field_type_7_is_repeated : _GEN_617; // @[Conditional.scala 39:67 Control.scala 57:36]
  wire  _GEN_969 = _T_19 ? classmeta_reg_desc_state_field_type_8_is_host : _GEN_618; // @[Conditional.scala 39:67 Control.scala 57:36]
  wire [15:0] _GEN_970 = _T_19 ? classmeta_reg_desc_state_field_type_8_sub_class_id : _GEN_619; // @[Conditional.scala 39:67 Control.scala 57:36]
  wire [4:0] _GEN_971 = _T_19 ? classmeta_reg_desc_state_field_type_8_field_type : _GEN_620; // @[Conditional.scala 39:67 Control.scala 57:36]
  wire  _GEN_972 = _T_19 ? classmeta_reg_desc_state_field_type_8_is_repeated : _GEN_621; // @[Conditional.scala 39:67 Control.scala 57:36]
  wire  _GEN_973 = _T_19 ? classmeta_reg_desc_state_field_type_9_is_host : _GEN_622; // @[Conditional.scala 39:67 Control.scala 57:36]
  wire [15:0] _GEN_974 = _T_19 ? classmeta_reg_desc_state_field_type_9_sub_class_id : _GEN_623; // @[Conditional.scala 39:67 Control.scala 57:36]
  wire [4:0] _GEN_975 = _T_19 ? classmeta_reg_desc_state_field_type_9_field_type : _GEN_624; // @[Conditional.scala 39:67 Control.scala 57:36]
  wire  _GEN_976 = _T_19 ? classmeta_reg_desc_state_field_type_9_is_repeated : _GEN_625; // @[Conditional.scala 39:67 Control.scala 57:36]
  wire  _GEN_977 = _T_19 ? classmeta_reg_desc_state_field_type_10_is_host : _GEN_626; // @[Conditional.scala 39:67 Control.scala 57:36]
  wire [15:0] _GEN_978 = _T_19 ? classmeta_reg_desc_state_field_type_10_sub_class_id : _GEN_627; // @[Conditional.scala 39:67 Control.scala 57:36]
  wire [4:0] _GEN_979 = _T_19 ? classmeta_reg_desc_state_field_type_10_field_type : _GEN_628; // @[Conditional.scala 39:67 Control.scala 57:36]
  wire  _GEN_980 = _T_19 ? classmeta_reg_desc_state_field_type_10_is_repeated : _GEN_629; // @[Conditional.scala 39:67 Control.scala 57:36]
  wire  _GEN_981 = _T_19 ? classmeta_reg_desc_state_field_type_11_is_host : _GEN_630; // @[Conditional.scala 39:67 Control.scala 57:36]
  wire [15:0] _GEN_982 = _T_19 ? classmeta_reg_desc_state_field_type_11_sub_class_id : _GEN_631; // @[Conditional.scala 39:67 Control.scala 57:36]
  wire [4:0] _GEN_983 = _T_19 ? classmeta_reg_desc_state_field_type_11_field_type : _GEN_632; // @[Conditional.scala 39:67 Control.scala 57:36]
  wire  _GEN_984 = _T_19 ? classmeta_reg_desc_state_field_type_11_is_repeated : _GEN_633; // @[Conditional.scala 39:67 Control.scala 57:36]
  wire  _GEN_985 = _T_19 ? classmeta_reg_desc_state_field_type_12_is_host : _GEN_634; // @[Conditional.scala 39:67 Control.scala 57:36]
  wire [15:0] _GEN_986 = _T_19 ? classmeta_reg_desc_state_field_type_12_sub_class_id : _GEN_635; // @[Conditional.scala 39:67 Control.scala 57:36]
  wire [4:0] _GEN_987 = _T_19 ? classmeta_reg_desc_state_field_type_12_field_type : _GEN_636; // @[Conditional.scala 39:67 Control.scala 57:36]
  wire  _GEN_988 = _T_19 ? classmeta_reg_desc_state_field_type_12_is_repeated : _GEN_637; // @[Conditional.scala 39:67 Control.scala 57:36]
  wire  _GEN_989 = _T_19 ? classmeta_reg_desc_state_field_type_13_is_host : _GEN_638; // @[Conditional.scala 39:67 Control.scala 57:36]
  wire [15:0] _GEN_990 = _T_19 ? classmeta_reg_desc_state_field_type_13_sub_class_id : _GEN_639; // @[Conditional.scala 39:67 Control.scala 57:36]
  wire [4:0] _GEN_991 = _T_19 ? classmeta_reg_desc_state_field_type_13_field_type : _GEN_640; // @[Conditional.scala 39:67 Control.scala 57:36]
  wire  _GEN_992 = _T_19 ? classmeta_reg_desc_state_field_type_13_is_repeated : _GEN_641; // @[Conditional.scala 39:67 Control.scala 57:36]
  wire [7:0] _GEN_1005 = _T_19 ? classmeta_reg_desc_state_max_field_num : _GEN_718; // @[Conditional.scala 39:67 Control.scala 57:36]
  wire [15:0] _GEN_1006 = _T_19 ? classmeta_reg_desc_state_class_length : _GEN_719; // @[Conditional.scala 39:67 Control.scala 57:36]
  wire [9:0] _GEN_1007 = _T_19 ? classmeta_reg_class_id : _GEN_720; // @[Conditional.scala 39:67 Control.scala 57:36]
  wire  _GEN_1008 = _T_19 ? 1'h0 : _GEN_722; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [10:0] _GEN_1009 = _T_19 ? 11'h0 : _GEN_723; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [63:0] _GEN_1010 = _T_19 ? 64'h0 : _GEN_724; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [10:0] _GEN_1022 = _T_17 ? _GEN_12 : {{1'd0}, _GEN_1007}; // @[Conditional.scala 39:67]
  wire [15:0] _GEN_1023 = _T_17 ? _GEN_13 : {{8'd0}, _GEN_1005}; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_1024 = _T_17 ? _GEN_14 : {{16'd0}, _GEN_1006}; // @[Conditional.scala 39:67]
  wire  _GEN_1146 = _T_17 ? 1'h0 : _GEN_801; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire  _GEN_1147 = _T_17 ? 1'h0 : _GEN_802; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [15:0] _GEN_1148 = _T_17 ? 16'h0 : _GEN_803; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [4:0] _GEN_1149 = _T_17 ? 5'h0 : _GEN_804; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire  _GEN_1150 = _T_17 ? 1'h0 : _GEN_805; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire  _GEN_1151 = _T_17 ? 1'h0 : _GEN_806; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [15:0] _GEN_1152 = _T_17 ? 16'h0 : _GEN_807; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [4:0] _GEN_1153 = _T_17 ? 5'h0 : _GEN_808; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire  _GEN_1154 = _T_17 ? 1'h0 : _GEN_809; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire  _GEN_1155 = _T_17 ? 1'h0 : _GEN_810; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [15:0] _GEN_1156 = _T_17 ? 16'h0 : _GEN_811; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [4:0] _GEN_1157 = _T_17 ? 5'h0 : _GEN_812; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire  _GEN_1158 = _T_17 ? 1'h0 : _GEN_813; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire  _GEN_1159 = _T_17 ? 1'h0 : _GEN_814; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [15:0] _GEN_1160 = _T_17 ? 16'h0 : _GEN_815; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [4:0] _GEN_1161 = _T_17 ? 5'h0 : _GEN_816; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire  _GEN_1162 = _T_17 ? 1'h0 : _GEN_817; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire  _GEN_1163 = _T_17 ? 1'h0 : _GEN_818; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [15:0] _GEN_1164 = _T_17 ? 16'h0 : _GEN_819; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [4:0] _GEN_1165 = _T_17 ? 5'h0 : _GEN_820; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire  _GEN_1166 = _T_17 ? 1'h0 : _GEN_821; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire  _GEN_1167 = _T_17 ? 1'h0 : _GEN_822; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [15:0] _GEN_1168 = _T_17 ? 16'h0 : _GEN_823; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [4:0] _GEN_1169 = _T_17 ? 5'h0 : _GEN_824; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire  _GEN_1170 = _T_17 ? 1'h0 : _GEN_825; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire  _GEN_1171 = _T_17 ? 1'h0 : _GEN_826; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [15:0] _GEN_1172 = _T_17 ? 16'h0 : _GEN_827; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [4:0] _GEN_1173 = _T_17 ? 5'h0 : _GEN_828; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire  _GEN_1174 = _T_17 ? 1'h0 : _GEN_829; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire  _GEN_1175 = _T_17 ? 1'h0 : _GEN_830; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [15:0] _GEN_1176 = _T_17 ? 16'h0 : _GEN_831; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [4:0] _GEN_1177 = _T_17 ? 5'h0 : _GEN_832; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire  _GEN_1178 = _T_17 ? 1'h0 : _GEN_833; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire  _GEN_1179 = _T_17 ? 1'h0 : _GEN_834; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [15:0] _GEN_1180 = _T_17 ? 16'h0 : _GEN_835; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [4:0] _GEN_1181 = _T_17 ? 5'h0 : _GEN_836; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire  _GEN_1182 = _T_17 ? 1'h0 : _GEN_837; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire  _GEN_1183 = _T_17 ? 1'h0 : _GEN_838; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [15:0] _GEN_1184 = _T_17 ? 16'h0 : _GEN_839; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [4:0] _GEN_1185 = _T_17 ? 5'h0 : _GEN_840; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire  _GEN_1186 = _T_17 ? 1'h0 : _GEN_841; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire  _GEN_1187 = _T_17 ? 1'h0 : _GEN_842; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [15:0] _GEN_1188 = _T_17 ? 16'h0 : _GEN_843; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [4:0] _GEN_1189 = _T_17 ? 5'h0 : _GEN_844; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire  _GEN_1190 = _T_17 ? 1'h0 : _GEN_845; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire  _GEN_1191 = _T_17 ? 1'h0 : _GEN_846; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [15:0] _GEN_1192 = _T_17 ? 16'h0 : _GEN_847; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [4:0] _GEN_1193 = _T_17 ? 5'h0 : _GEN_848; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire  _GEN_1194 = _T_17 ? 1'h0 : _GEN_849; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire  _GEN_1195 = _T_17 ? 1'h0 : _GEN_850; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [15:0] _GEN_1196 = _T_17 ? 16'h0 : _GEN_851; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [4:0] _GEN_1197 = _T_17 ? 5'h0 : _GEN_852; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire  _GEN_1198 = _T_17 ? 1'h0 : _GEN_853; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire  _GEN_1199 = _T_17 ? 1'h0 : _GEN_854; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [15:0] _GEN_1200 = _T_17 ? 16'h0 : _GEN_855; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [4:0] _GEN_1201 = _T_17 ? 5'h0 : _GEN_856; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire  _GEN_1202 = _T_17 ? 1'h0 : _GEN_857; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire  _GEN_1203 = _T_17 ? 1'h0 : _GEN_858; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [15:0] _GEN_1204 = _T_17 ? 16'h0 : _GEN_859; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [4:0] _GEN_1205 = _T_17 ? 5'h0 : _GEN_860; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire  _GEN_1206 = _T_17 ? 1'h0 : _GEN_861; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire  _GEN_1207 = _T_17 ? 1'h0 : _GEN_862; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [15:0] _GEN_1208 = _T_17 ? 16'h0 : _GEN_863; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [4:0] _GEN_1209 = _T_17 ? 5'h0 : _GEN_864; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire  _GEN_1210 = _T_17 ? 1'h0 : _GEN_865; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire  _GEN_1211 = _T_17 ? 1'h0 : _GEN_866; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [15:0] _GEN_1212 = _T_17 ? 16'h0 : _GEN_867; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [4:0] _GEN_1213 = _T_17 ? 5'h0 : _GEN_868; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire  _GEN_1214 = _T_17 ? 1'h0 : _GEN_869; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire  _GEN_1215 = _T_17 ? 1'h0 : _GEN_870; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [15:0] _GEN_1216 = _T_17 ? 16'h0 : _GEN_871; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [4:0] _GEN_1217 = _T_17 ? 5'h0 : _GEN_872; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire  _GEN_1218 = _T_17 ? 1'h0 : _GEN_873; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire  _GEN_1219 = _T_17 ? 1'h0 : _GEN_874; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [15:0] _GEN_1220 = _T_17 ? 16'h0 : _GEN_875; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [4:0] _GEN_1221 = _T_17 ? 5'h0 : _GEN_876; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire  _GEN_1222 = _T_17 ? 1'h0 : _GEN_877; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire  _GEN_1223 = _T_17 ? 1'h0 : _GEN_878; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [15:0] _GEN_1224 = _T_17 ? 16'h0 : _GEN_879; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [4:0] _GEN_1225 = _T_17 ? 5'h0 : _GEN_880; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire  _GEN_1226 = _T_17 ? 1'h0 : _GEN_881; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire  _GEN_1227 = _T_17 ? 1'h0 : _GEN_882; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [15:0] _GEN_1228 = _T_17 ? 16'h0 : _GEN_883; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [4:0] _GEN_1229 = _T_17 ? 5'h0 : _GEN_884; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire  _GEN_1230 = _T_17 ? 1'h0 : _GEN_885; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire  _GEN_1231 = _T_17 ? 1'h0 : _GEN_886; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [15:0] _GEN_1232 = _T_17 ? 16'h0 : _GEN_887; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [4:0] _GEN_1233 = _T_17 ? 5'h0 : _GEN_888; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire  _GEN_1234 = _T_17 ? 1'h0 : _GEN_889; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire  _GEN_1235 = _T_17 ? 1'h0 : _GEN_890; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [15:0] _GEN_1236 = _T_17 ? 16'h0 : _GEN_891; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [4:0] _GEN_1237 = _T_17 ? 5'h0 : _GEN_892; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire  _GEN_1238 = _T_17 ? 1'h0 : _GEN_893; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire  _GEN_1239 = _T_17 ? 1'h0 : _GEN_894; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [15:0] _GEN_1240 = _T_17 ? 16'h0 : _GEN_895; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [4:0] _GEN_1241 = _T_17 ? 5'h0 : _GEN_896; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire  _GEN_1242 = _T_17 ? 1'h0 : _GEN_897; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire  _GEN_1243 = _T_17 ? 1'h0 : _GEN_898; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [15:0] _GEN_1244 = _T_17 ? 16'h0 : _GEN_899; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [4:0] _GEN_1245 = _T_17 ? 5'h0 : _GEN_900; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire  _GEN_1246 = _T_17 ? 1'h0 : _GEN_901; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire  _GEN_1247 = _T_17 ? 1'h0 : _GEN_902; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [15:0] _GEN_1248 = _T_17 ? 16'h0 : _GEN_903; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [4:0] _GEN_1249 = _T_17 ? 5'h0 : _GEN_904; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire  _GEN_1250 = _T_17 ? 1'h0 : _GEN_905; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire  _GEN_1251 = _T_17 ? 1'h0 : _GEN_906; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [15:0] _GEN_1252 = _T_17 ? 16'h0 : _GEN_907; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [4:0] _GEN_1253 = _T_17 ? 5'h0 : _GEN_908; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire  _GEN_1254 = _T_17 ? 1'h0 : _GEN_909; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire  _GEN_1255 = _T_17 ? 1'h0 : _GEN_910; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [15:0] _GEN_1256 = _T_17 ? 16'h0 : _GEN_911; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [4:0] _GEN_1257 = _T_17 ? 5'h0 : _GEN_912; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire  _GEN_1258 = _T_17 ? 1'h0 : _GEN_913; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire  _GEN_1259 = _T_17 ? 1'h0 : _GEN_914; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [15:0] _GEN_1260 = _T_17 ? 16'h0 : _GEN_915; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [4:0] _GEN_1261 = _T_17 ? 5'h0 : _GEN_916; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire  _GEN_1262 = _T_17 ? 1'h0 : _GEN_917; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire  _GEN_1263 = _T_17 ? 1'h0 : _GEN_918; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [15:0] _GEN_1264 = _T_17 ? 16'h0 : _GEN_919; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [4:0] _GEN_1265 = _T_17 ? 5'h0 : _GEN_920; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire  _GEN_1266 = _T_17 ? 1'h0 : _GEN_921; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire  _GEN_1267 = _T_17 ? 1'h0 : _GEN_922; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [15:0] _GEN_1268 = _T_17 ? 16'h0 : _GEN_923; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [4:0] _GEN_1269 = _T_17 ? 5'h0 : _GEN_924; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire  _GEN_1270 = _T_17 ? 1'h0 : _GEN_925; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire  _GEN_1271 = _T_17 ? 1'h0 : _GEN_926; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [15:0] _GEN_1272 = _T_17 ? 16'h0 : _GEN_927; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [4:0] _GEN_1273 = _T_17 ? 5'h0 : _GEN_928; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire  _GEN_1274 = _T_17 ? 1'h0 : _GEN_929; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire  _GEN_1275 = _T_17 ? 1'h0 : _GEN_930; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [15:0] _GEN_1276 = _T_17 ? 16'h0 : _GEN_931; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [4:0] _GEN_1277 = _T_17 ? 5'h0 : _GEN_932; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire  _GEN_1278 = _T_17 ? 1'h0 : _GEN_933; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [7:0] _GEN_1279 = _T_17 ? 8'h0 : _GEN_934; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [15:0] _GEN_1280 = _T_17 ? 16'h0 : _GEN_935; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [9:0] _GEN_1281 = _T_17 ? 10'h0 : _GEN_936; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire  _GEN_1294 = _T_17 ? 1'h0 : _GEN_1008; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [10:0] _GEN_1295 = _T_17 ? 11'h0 : _GEN_1009; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [63:0] _GEN_1296 = _T_17 ? 64'h0 : _GEN_1010; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [10:0] _GEN_1311 = _T_15 ? {{1'd0}, classmeta_reg_class_id} : _GEN_1022; // @[Conditional.scala 39:67 Control.scala 57:36]
  wire [15:0] _GEN_1312 = _T_15 ? {{8'd0}, classmeta_reg_desc_state_max_field_num} : _GEN_1023; // @[Conditional.scala 39:67 Control.scala 57:36]
  wire [31:0] _GEN_1313 = _T_15 ? {{16'd0}, classmeta_reg_desc_state_class_length} : _GEN_1024; // @[Conditional.scala 39:67 Control.scala 57:36]
  wire  _GEN_1434 = _T_15 ? 1'h0 : _GEN_1146; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire  _GEN_1435 = _T_15 ? 1'h0 : _GEN_1147; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [15:0] _GEN_1436 = _T_15 ? 16'h0 : _GEN_1148; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [4:0] _GEN_1437 = _T_15 ? 5'h0 : _GEN_1149; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire  _GEN_1438 = _T_15 ? 1'h0 : _GEN_1150; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire  _GEN_1439 = _T_15 ? 1'h0 : _GEN_1151; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [15:0] _GEN_1440 = _T_15 ? 16'h0 : _GEN_1152; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [4:0] _GEN_1441 = _T_15 ? 5'h0 : _GEN_1153; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire  _GEN_1442 = _T_15 ? 1'h0 : _GEN_1154; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire  _GEN_1443 = _T_15 ? 1'h0 : _GEN_1155; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [15:0] _GEN_1444 = _T_15 ? 16'h0 : _GEN_1156; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [4:0] _GEN_1445 = _T_15 ? 5'h0 : _GEN_1157; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire  _GEN_1446 = _T_15 ? 1'h0 : _GEN_1158; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire  _GEN_1447 = _T_15 ? 1'h0 : _GEN_1159; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [15:0] _GEN_1448 = _T_15 ? 16'h0 : _GEN_1160; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [4:0] _GEN_1449 = _T_15 ? 5'h0 : _GEN_1161; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire  _GEN_1450 = _T_15 ? 1'h0 : _GEN_1162; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire  _GEN_1451 = _T_15 ? 1'h0 : _GEN_1163; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [15:0] _GEN_1452 = _T_15 ? 16'h0 : _GEN_1164; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [4:0] _GEN_1453 = _T_15 ? 5'h0 : _GEN_1165; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire  _GEN_1454 = _T_15 ? 1'h0 : _GEN_1166; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire  _GEN_1455 = _T_15 ? 1'h0 : _GEN_1167; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [15:0] _GEN_1456 = _T_15 ? 16'h0 : _GEN_1168; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [4:0] _GEN_1457 = _T_15 ? 5'h0 : _GEN_1169; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire  _GEN_1458 = _T_15 ? 1'h0 : _GEN_1170; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire  _GEN_1459 = _T_15 ? 1'h0 : _GEN_1171; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [15:0] _GEN_1460 = _T_15 ? 16'h0 : _GEN_1172; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [4:0] _GEN_1461 = _T_15 ? 5'h0 : _GEN_1173; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire  _GEN_1462 = _T_15 ? 1'h0 : _GEN_1174; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire  _GEN_1463 = _T_15 ? 1'h0 : _GEN_1175; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [15:0] _GEN_1464 = _T_15 ? 16'h0 : _GEN_1176; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [4:0] _GEN_1465 = _T_15 ? 5'h0 : _GEN_1177; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire  _GEN_1466 = _T_15 ? 1'h0 : _GEN_1178; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire  _GEN_1467 = _T_15 ? 1'h0 : _GEN_1179; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [15:0] _GEN_1468 = _T_15 ? 16'h0 : _GEN_1180; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [4:0] _GEN_1469 = _T_15 ? 5'h0 : _GEN_1181; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire  _GEN_1470 = _T_15 ? 1'h0 : _GEN_1182; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire  _GEN_1471 = _T_15 ? 1'h0 : _GEN_1183; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [15:0] _GEN_1472 = _T_15 ? 16'h0 : _GEN_1184; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [4:0] _GEN_1473 = _T_15 ? 5'h0 : _GEN_1185; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire  _GEN_1474 = _T_15 ? 1'h0 : _GEN_1186; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire  _GEN_1475 = _T_15 ? 1'h0 : _GEN_1187; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [15:0] _GEN_1476 = _T_15 ? 16'h0 : _GEN_1188; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [4:0] _GEN_1477 = _T_15 ? 5'h0 : _GEN_1189; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire  _GEN_1478 = _T_15 ? 1'h0 : _GEN_1190; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire  _GEN_1479 = _T_15 ? 1'h0 : _GEN_1191; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [15:0] _GEN_1480 = _T_15 ? 16'h0 : _GEN_1192; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [4:0] _GEN_1481 = _T_15 ? 5'h0 : _GEN_1193; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire  _GEN_1482 = _T_15 ? 1'h0 : _GEN_1194; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire  _GEN_1483 = _T_15 ? 1'h0 : _GEN_1195; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [15:0] _GEN_1484 = _T_15 ? 16'h0 : _GEN_1196; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [4:0] _GEN_1485 = _T_15 ? 5'h0 : _GEN_1197; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire  _GEN_1486 = _T_15 ? 1'h0 : _GEN_1198; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire  _GEN_1487 = _T_15 ? 1'h0 : _GEN_1199; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [15:0] _GEN_1488 = _T_15 ? 16'h0 : _GEN_1200; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [4:0] _GEN_1489 = _T_15 ? 5'h0 : _GEN_1201; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire  _GEN_1490 = _T_15 ? 1'h0 : _GEN_1202; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire  _GEN_1491 = _T_15 ? 1'h0 : _GEN_1203; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [15:0] _GEN_1492 = _T_15 ? 16'h0 : _GEN_1204; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [4:0] _GEN_1493 = _T_15 ? 5'h0 : _GEN_1205; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire  _GEN_1494 = _T_15 ? 1'h0 : _GEN_1206; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire  _GEN_1495 = _T_15 ? 1'h0 : _GEN_1207; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [15:0] _GEN_1496 = _T_15 ? 16'h0 : _GEN_1208; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [4:0] _GEN_1497 = _T_15 ? 5'h0 : _GEN_1209; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire  _GEN_1498 = _T_15 ? 1'h0 : _GEN_1210; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire  _GEN_1499 = _T_15 ? 1'h0 : _GEN_1211; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [15:0] _GEN_1500 = _T_15 ? 16'h0 : _GEN_1212; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [4:0] _GEN_1501 = _T_15 ? 5'h0 : _GEN_1213; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire  _GEN_1502 = _T_15 ? 1'h0 : _GEN_1214; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire  _GEN_1503 = _T_15 ? 1'h0 : _GEN_1215; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [15:0] _GEN_1504 = _T_15 ? 16'h0 : _GEN_1216; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [4:0] _GEN_1505 = _T_15 ? 5'h0 : _GEN_1217; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire  _GEN_1506 = _T_15 ? 1'h0 : _GEN_1218; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire  _GEN_1507 = _T_15 ? 1'h0 : _GEN_1219; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [15:0] _GEN_1508 = _T_15 ? 16'h0 : _GEN_1220; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [4:0] _GEN_1509 = _T_15 ? 5'h0 : _GEN_1221; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire  _GEN_1510 = _T_15 ? 1'h0 : _GEN_1222; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire  _GEN_1511 = _T_15 ? 1'h0 : _GEN_1223; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [15:0] _GEN_1512 = _T_15 ? 16'h0 : _GEN_1224; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [4:0] _GEN_1513 = _T_15 ? 5'h0 : _GEN_1225; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire  _GEN_1514 = _T_15 ? 1'h0 : _GEN_1226; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire  _GEN_1515 = _T_15 ? 1'h0 : _GEN_1227; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [15:0] _GEN_1516 = _T_15 ? 16'h0 : _GEN_1228; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [4:0] _GEN_1517 = _T_15 ? 5'h0 : _GEN_1229; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire  _GEN_1518 = _T_15 ? 1'h0 : _GEN_1230; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire  _GEN_1519 = _T_15 ? 1'h0 : _GEN_1231; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [15:0] _GEN_1520 = _T_15 ? 16'h0 : _GEN_1232; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [4:0] _GEN_1521 = _T_15 ? 5'h0 : _GEN_1233; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire  _GEN_1522 = _T_15 ? 1'h0 : _GEN_1234; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire  _GEN_1523 = _T_15 ? 1'h0 : _GEN_1235; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [15:0] _GEN_1524 = _T_15 ? 16'h0 : _GEN_1236; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [4:0] _GEN_1525 = _T_15 ? 5'h0 : _GEN_1237; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire  _GEN_1526 = _T_15 ? 1'h0 : _GEN_1238; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire  _GEN_1527 = _T_15 ? 1'h0 : _GEN_1239; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [15:0] _GEN_1528 = _T_15 ? 16'h0 : _GEN_1240; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [4:0] _GEN_1529 = _T_15 ? 5'h0 : _GEN_1241; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire  _GEN_1530 = _T_15 ? 1'h0 : _GEN_1242; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire  _GEN_1531 = _T_15 ? 1'h0 : _GEN_1243; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [15:0] _GEN_1532 = _T_15 ? 16'h0 : _GEN_1244; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [4:0] _GEN_1533 = _T_15 ? 5'h0 : _GEN_1245; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire  _GEN_1534 = _T_15 ? 1'h0 : _GEN_1246; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire  _GEN_1535 = _T_15 ? 1'h0 : _GEN_1247; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [15:0] _GEN_1536 = _T_15 ? 16'h0 : _GEN_1248; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [4:0] _GEN_1537 = _T_15 ? 5'h0 : _GEN_1249; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire  _GEN_1538 = _T_15 ? 1'h0 : _GEN_1250; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire  _GEN_1539 = _T_15 ? 1'h0 : _GEN_1251; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [15:0] _GEN_1540 = _T_15 ? 16'h0 : _GEN_1252; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [4:0] _GEN_1541 = _T_15 ? 5'h0 : _GEN_1253; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire  _GEN_1542 = _T_15 ? 1'h0 : _GEN_1254; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire  _GEN_1543 = _T_15 ? 1'h0 : _GEN_1255; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [15:0] _GEN_1544 = _T_15 ? 16'h0 : _GEN_1256; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [4:0] _GEN_1545 = _T_15 ? 5'h0 : _GEN_1257; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire  _GEN_1546 = _T_15 ? 1'h0 : _GEN_1258; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire  _GEN_1547 = _T_15 ? 1'h0 : _GEN_1259; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [15:0] _GEN_1548 = _T_15 ? 16'h0 : _GEN_1260; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [4:0] _GEN_1549 = _T_15 ? 5'h0 : _GEN_1261; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire  _GEN_1550 = _T_15 ? 1'h0 : _GEN_1262; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire  _GEN_1551 = _T_15 ? 1'h0 : _GEN_1263; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [15:0] _GEN_1552 = _T_15 ? 16'h0 : _GEN_1264; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [4:0] _GEN_1553 = _T_15 ? 5'h0 : _GEN_1265; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire  _GEN_1554 = _T_15 ? 1'h0 : _GEN_1266; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire  _GEN_1555 = _T_15 ? 1'h0 : _GEN_1267; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [15:0] _GEN_1556 = _T_15 ? 16'h0 : _GEN_1268; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [4:0] _GEN_1557 = _T_15 ? 5'h0 : _GEN_1269; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire  _GEN_1558 = _T_15 ? 1'h0 : _GEN_1270; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire  _GEN_1559 = _T_15 ? 1'h0 : _GEN_1271; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [15:0] _GEN_1560 = _T_15 ? 16'h0 : _GEN_1272; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [4:0] _GEN_1561 = _T_15 ? 5'h0 : _GEN_1273; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire  _GEN_1562 = _T_15 ? 1'h0 : _GEN_1274; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire  _GEN_1563 = _T_15 ? 1'h0 : _GEN_1275; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [15:0] _GEN_1564 = _T_15 ? 16'h0 : _GEN_1276; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [4:0] _GEN_1565 = _T_15 ? 5'h0 : _GEN_1277; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire  _GEN_1566 = _T_15 ? 1'h0 : _GEN_1278; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [7:0] _GEN_1567 = _T_15 ? 8'h0 : _GEN_1279; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [15:0] _GEN_1568 = _T_15 ? 16'h0 : _GEN_1280; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [9:0] _GEN_1569 = _T_15 ? 10'h0 : _GEN_1281; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire  _GEN_1582 = _T_15 ? 1'h0 : _GEN_1294; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [10:0] _GEN_1583 = _T_15 ? 11'h0 : _GEN_1295; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [63:0] _GEN_1584 = _T_15 ? 64'h0 : _GEN_1296; // @[Conditional.scala 39:67 Util.scala 13:25]
  wire [10:0] _GEN_1600 = _T_1 ? {{1'd0}, classmeta_reg_class_id} : _GEN_1311; // @[Conditional.scala 40:58 Control.scala 57:36]
  wire [15:0] _GEN_1601 = _T_1 ? {{8'd0}, classmeta_reg_desc_state_max_field_num} : _GEN_1312; // @[Conditional.scala 40:58 Control.scala 57:36]
  wire [31:0] _GEN_1602 = _T_1 ? {{16'd0}, classmeta_reg_desc_state_class_length} : _GEN_1313; // @[Conditional.scala 40:58 Control.scala 57:36]
  wire [10:0] _GEN_1872 = _T_1 ? 11'h0 : _GEN_1583; // @[Conditional.scala 40:58 Util.scala 13:25]
  assign io_axi_aw_ready = s_wr == 3'h0; // @[Control.scala 69:34]
  assign io_axi_w_ready = s_wr == 3'h1 | s_wr == 3'h2 | s_wr == 3'h3 | s_wr == 3'h4 | s_wr == 3'h5 | s_wr == 3'h6 &
    io_ser_cmd_ready | s_wr == 3'h7; // @[Control.scala 70:244]
  assign io_axi_r_valid = 1'h1; // @[Control.scala 64:25]
  assign io_axi_r_bits_data = {{480'd0}, cur_data}; // @[Control.scala 65:25]
  assign io_metadata_init_valid = _T_1 ? 1'h0 : _GEN_1434; // @[Conditional.scala 40:58 Util.scala 13:25]
  assign io_metadata_init_bits_class_id = _T_1 ? 10'h0 : _GEN_1569; // @[Conditional.scala 40:58 Util.scala 13:25]
  assign io_metadata_init_bits_desc_state_class_length = _T_1 ? 16'h0 : _GEN_1568; // @[Conditional.scala 40:58 Util.scala 13:25]
  assign io_metadata_init_bits_desc_state_max_field_num = _T_1 ? 8'h0 : _GEN_1567; // @[Conditional.scala 40:58 Util.scala 13:25]
  assign io_metadata_init_bits_desc_state_field_type_0_is_repeated = _T_1 ? 1'h0 : _GEN_1438; // @[Conditional.scala 40:58 Util.scala 13:25]
  assign io_metadata_init_bits_desc_state_field_type_0_field_type = _T_1 ? 5'h0 : _GEN_1437; // @[Conditional.scala 40:58 Util.scala 13:25]
  assign io_metadata_init_bits_desc_state_field_type_0_sub_class_id = _T_1 ? 16'h0 : _GEN_1436; // @[Conditional.scala 40:58 Util.scala 13:25]
  assign io_metadata_init_bits_desc_state_field_type_0_is_host = _T_1 ? 1'h0 : _GEN_1435; // @[Conditional.scala 40:58 Util.scala 13:25]
  assign io_metadata_init_bits_desc_state_field_type_1_is_repeated = _T_1 ? 1'h0 : _GEN_1442; // @[Conditional.scala 40:58 Util.scala 13:25]
  assign io_metadata_init_bits_desc_state_field_type_1_field_type = _T_1 ? 5'h0 : _GEN_1441; // @[Conditional.scala 40:58 Util.scala 13:25]
  assign io_metadata_init_bits_desc_state_field_type_1_sub_class_id = _T_1 ? 16'h0 : _GEN_1440; // @[Conditional.scala 40:58 Util.scala 13:25]
  assign io_metadata_init_bits_desc_state_field_type_1_is_host = _T_1 ? 1'h0 : _GEN_1439; // @[Conditional.scala 40:58 Util.scala 13:25]
  assign io_metadata_init_bits_desc_state_field_type_2_is_repeated = _T_1 ? 1'h0 : _GEN_1446; // @[Conditional.scala 40:58 Util.scala 13:25]
  assign io_metadata_init_bits_desc_state_field_type_2_field_type = _T_1 ? 5'h0 : _GEN_1445; // @[Conditional.scala 40:58 Util.scala 13:25]
  assign io_metadata_init_bits_desc_state_field_type_2_sub_class_id = _T_1 ? 16'h0 : _GEN_1444; // @[Conditional.scala 40:58 Util.scala 13:25]
  assign io_metadata_init_bits_desc_state_field_type_2_is_host = _T_1 ? 1'h0 : _GEN_1443; // @[Conditional.scala 40:58 Util.scala 13:25]
  assign io_metadata_init_bits_desc_state_field_type_3_is_repeated = _T_1 ? 1'h0 : _GEN_1450; // @[Conditional.scala 40:58 Util.scala 13:25]
  assign io_metadata_init_bits_desc_state_field_type_3_field_type = _T_1 ? 5'h0 : _GEN_1449; // @[Conditional.scala 40:58 Util.scala 13:25]
  assign io_metadata_init_bits_desc_state_field_type_3_sub_class_id = _T_1 ? 16'h0 : _GEN_1448; // @[Conditional.scala 40:58 Util.scala 13:25]
  assign io_metadata_init_bits_desc_state_field_type_3_is_host = _T_1 ? 1'h0 : _GEN_1447; // @[Conditional.scala 40:58 Util.scala 13:25]
  assign io_metadata_init_bits_desc_state_field_type_4_is_repeated = _T_1 ? 1'h0 : _GEN_1454; // @[Conditional.scala 40:58 Util.scala 13:25]
  assign io_metadata_init_bits_desc_state_field_type_4_field_type = _T_1 ? 5'h0 : _GEN_1453; // @[Conditional.scala 40:58 Util.scala 13:25]
  assign io_metadata_init_bits_desc_state_field_type_4_sub_class_id = _T_1 ? 16'h0 : _GEN_1452; // @[Conditional.scala 40:58 Util.scala 13:25]
  assign io_metadata_init_bits_desc_state_field_type_4_is_host = _T_1 ? 1'h0 : _GEN_1451; // @[Conditional.scala 40:58 Util.scala 13:25]
  assign io_metadata_init_bits_desc_state_field_type_5_is_repeated = _T_1 ? 1'h0 : _GEN_1458; // @[Conditional.scala 40:58 Util.scala 13:25]
  assign io_metadata_init_bits_desc_state_field_type_5_field_type = _T_1 ? 5'h0 : _GEN_1457; // @[Conditional.scala 40:58 Util.scala 13:25]
  assign io_metadata_init_bits_desc_state_field_type_5_sub_class_id = _T_1 ? 16'h0 : _GEN_1456; // @[Conditional.scala 40:58 Util.scala 13:25]
  assign io_metadata_init_bits_desc_state_field_type_5_is_host = _T_1 ? 1'h0 : _GEN_1455; // @[Conditional.scala 40:58 Util.scala 13:25]
  assign io_metadata_init_bits_desc_state_field_type_6_is_repeated = _T_1 ? 1'h0 : _GEN_1462; // @[Conditional.scala 40:58 Util.scala 13:25]
  assign io_metadata_init_bits_desc_state_field_type_6_field_type = _T_1 ? 5'h0 : _GEN_1461; // @[Conditional.scala 40:58 Util.scala 13:25]
  assign io_metadata_init_bits_desc_state_field_type_6_sub_class_id = _T_1 ? 16'h0 : _GEN_1460; // @[Conditional.scala 40:58 Util.scala 13:25]
  assign io_metadata_init_bits_desc_state_field_type_6_is_host = _T_1 ? 1'h0 : _GEN_1459; // @[Conditional.scala 40:58 Util.scala 13:25]
  assign io_metadata_init_bits_desc_state_field_type_7_is_repeated = _T_1 ? 1'h0 : _GEN_1466; // @[Conditional.scala 40:58 Util.scala 13:25]
  assign io_metadata_init_bits_desc_state_field_type_7_field_type = _T_1 ? 5'h0 : _GEN_1465; // @[Conditional.scala 40:58 Util.scala 13:25]
  assign io_metadata_init_bits_desc_state_field_type_7_sub_class_id = _T_1 ? 16'h0 : _GEN_1464; // @[Conditional.scala 40:58 Util.scala 13:25]
  assign io_metadata_init_bits_desc_state_field_type_7_is_host = _T_1 ? 1'h0 : _GEN_1463; // @[Conditional.scala 40:58 Util.scala 13:25]
  assign io_metadata_init_bits_desc_state_field_type_8_is_repeated = _T_1 ? 1'h0 : _GEN_1470; // @[Conditional.scala 40:58 Util.scala 13:25]
  assign io_metadata_init_bits_desc_state_field_type_8_field_type = _T_1 ? 5'h0 : _GEN_1469; // @[Conditional.scala 40:58 Util.scala 13:25]
  assign io_metadata_init_bits_desc_state_field_type_8_sub_class_id = _T_1 ? 16'h0 : _GEN_1468; // @[Conditional.scala 40:58 Util.scala 13:25]
  assign io_metadata_init_bits_desc_state_field_type_8_is_host = _T_1 ? 1'h0 : _GEN_1467; // @[Conditional.scala 40:58 Util.scala 13:25]
  assign io_metadata_init_bits_desc_state_field_type_9_is_repeated = _T_1 ? 1'h0 : _GEN_1474; // @[Conditional.scala 40:58 Util.scala 13:25]
  assign io_metadata_init_bits_desc_state_field_type_9_field_type = _T_1 ? 5'h0 : _GEN_1473; // @[Conditional.scala 40:58 Util.scala 13:25]
  assign io_metadata_init_bits_desc_state_field_type_9_sub_class_id = _T_1 ? 16'h0 : _GEN_1472; // @[Conditional.scala 40:58 Util.scala 13:25]
  assign io_metadata_init_bits_desc_state_field_type_9_is_host = _T_1 ? 1'h0 : _GEN_1471; // @[Conditional.scala 40:58 Util.scala 13:25]
  assign io_metadata_init_bits_desc_state_field_type_10_is_repeated = _T_1 ? 1'h0 : _GEN_1478; // @[Conditional.scala 40:58 Util.scala 13:25]
  assign io_metadata_init_bits_desc_state_field_type_10_field_type = _T_1 ? 5'h0 : _GEN_1477; // @[Conditional.scala 40:58 Util.scala 13:25]
  assign io_metadata_init_bits_desc_state_field_type_10_sub_class_id = _T_1 ? 16'h0 : _GEN_1476; // @[Conditional.scala 40:58 Util.scala 13:25]
  assign io_metadata_init_bits_desc_state_field_type_10_is_host = _T_1 ? 1'h0 : _GEN_1475; // @[Conditional.scala 40:58 Util.scala 13:25]
  assign io_metadata_init_bits_desc_state_field_type_11_is_repeated = _T_1 ? 1'h0 : _GEN_1482; // @[Conditional.scala 40:58 Util.scala 13:25]
  assign io_metadata_init_bits_desc_state_field_type_11_field_type = _T_1 ? 5'h0 : _GEN_1481; // @[Conditional.scala 40:58 Util.scala 13:25]
  assign io_metadata_init_bits_desc_state_field_type_11_sub_class_id = _T_1 ? 16'h0 : _GEN_1480; // @[Conditional.scala 40:58 Util.scala 13:25]
  assign io_metadata_init_bits_desc_state_field_type_11_is_host = _T_1 ? 1'h0 : _GEN_1479; // @[Conditional.scala 40:58 Util.scala 13:25]
  assign io_metadata_init_bits_desc_state_field_type_12_is_repeated = _T_1 ? 1'h0 : _GEN_1486; // @[Conditional.scala 40:58 Util.scala 13:25]
  assign io_metadata_init_bits_desc_state_field_type_12_field_type = _T_1 ? 5'h0 : _GEN_1485; // @[Conditional.scala 40:58 Util.scala 13:25]
  assign io_metadata_init_bits_desc_state_field_type_12_sub_class_id = _T_1 ? 16'h0 : _GEN_1484; // @[Conditional.scala 40:58 Util.scala 13:25]
  assign io_metadata_init_bits_desc_state_field_type_12_is_host = _T_1 ? 1'h0 : _GEN_1483; // @[Conditional.scala 40:58 Util.scala 13:25]
  assign io_metadata_init_bits_desc_state_field_type_13_is_repeated = _T_1 ? 1'h0 : _GEN_1490; // @[Conditional.scala 40:58 Util.scala 13:25]
  assign io_metadata_init_bits_desc_state_field_type_13_field_type = _T_1 ? 5'h0 : _GEN_1489; // @[Conditional.scala 40:58 Util.scala 13:25]
  assign io_metadata_init_bits_desc_state_field_type_13_sub_class_id = _T_1 ? 16'h0 : _GEN_1488; // @[Conditional.scala 40:58 Util.scala 13:25]
  assign io_metadata_init_bits_desc_state_field_type_13_is_host = _T_1 ? 1'h0 : _GEN_1487; // @[Conditional.scala 40:58 Util.scala 13:25]
  assign io_metadata_init_bits_desc_state_field_type_14_is_repeated = _T_1 ? 1'h0 : _GEN_1494; // @[Conditional.scala 40:58 Util.scala 13:25]
  assign io_metadata_init_bits_desc_state_field_type_14_field_type = _T_1 ? 5'h0 : _GEN_1493; // @[Conditional.scala 40:58 Util.scala 13:25]
  assign io_metadata_init_bits_desc_state_field_type_14_sub_class_id = _T_1 ? 16'h0 : _GEN_1492; // @[Conditional.scala 40:58 Util.scala 13:25]
  assign io_metadata_init_bits_desc_state_field_type_14_is_host = _T_1 ? 1'h0 : _GEN_1491; // @[Conditional.scala 40:58 Util.scala 13:25]
  assign io_metadata_init_bits_desc_state_field_type_15_is_repeated = _T_1 ? 1'h0 : _GEN_1498; // @[Conditional.scala 40:58 Util.scala 13:25]
  assign io_metadata_init_bits_desc_state_field_type_15_field_type = _T_1 ? 5'h0 : _GEN_1497; // @[Conditional.scala 40:58 Util.scala 13:25]
  assign io_metadata_init_bits_desc_state_field_type_15_sub_class_id = _T_1 ? 16'h0 : _GEN_1496; // @[Conditional.scala 40:58 Util.scala 13:25]
  assign io_metadata_init_bits_desc_state_field_type_15_is_host = _T_1 ? 1'h0 : _GEN_1495; // @[Conditional.scala 40:58 Util.scala 13:25]
  assign io_metadata_init_bits_desc_state_field_type_16_is_repeated = _T_1 ? 1'h0 : _GEN_1502; // @[Conditional.scala 40:58 Util.scala 13:25]
  assign io_metadata_init_bits_desc_state_field_type_16_field_type = _T_1 ? 5'h0 : _GEN_1501; // @[Conditional.scala 40:58 Util.scala 13:25]
  assign io_metadata_init_bits_desc_state_field_type_16_sub_class_id = _T_1 ? 16'h0 : _GEN_1500; // @[Conditional.scala 40:58 Util.scala 13:25]
  assign io_metadata_init_bits_desc_state_field_type_16_is_host = _T_1 ? 1'h0 : _GEN_1499; // @[Conditional.scala 40:58 Util.scala 13:25]
  assign io_metadata_init_bits_desc_state_field_type_17_is_repeated = _T_1 ? 1'h0 : _GEN_1506; // @[Conditional.scala 40:58 Util.scala 13:25]
  assign io_metadata_init_bits_desc_state_field_type_17_field_type = _T_1 ? 5'h0 : _GEN_1505; // @[Conditional.scala 40:58 Util.scala 13:25]
  assign io_metadata_init_bits_desc_state_field_type_17_sub_class_id = _T_1 ? 16'h0 : _GEN_1504; // @[Conditional.scala 40:58 Util.scala 13:25]
  assign io_metadata_init_bits_desc_state_field_type_17_is_host = _T_1 ? 1'h0 : _GEN_1503; // @[Conditional.scala 40:58 Util.scala 13:25]
  assign io_metadata_init_bits_desc_state_field_type_18_is_repeated = _T_1 ? 1'h0 : _GEN_1510; // @[Conditional.scala 40:58 Util.scala 13:25]
  assign io_metadata_init_bits_desc_state_field_type_18_field_type = _T_1 ? 5'h0 : _GEN_1509; // @[Conditional.scala 40:58 Util.scala 13:25]
  assign io_metadata_init_bits_desc_state_field_type_18_sub_class_id = _T_1 ? 16'h0 : _GEN_1508; // @[Conditional.scala 40:58 Util.scala 13:25]
  assign io_metadata_init_bits_desc_state_field_type_18_is_host = _T_1 ? 1'h0 : _GEN_1507; // @[Conditional.scala 40:58 Util.scala 13:25]
  assign io_metadata_init_bits_desc_state_field_type_19_is_repeated = _T_1 ? 1'h0 : _GEN_1514; // @[Conditional.scala 40:58 Util.scala 13:25]
  assign io_metadata_init_bits_desc_state_field_type_19_field_type = _T_1 ? 5'h0 : _GEN_1513; // @[Conditional.scala 40:58 Util.scala 13:25]
  assign io_metadata_init_bits_desc_state_field_type_19_sub_class_id = _T_1 ? 16'h0 : _GEN_1512; // @[Conditional.scala 40:58 Util.scala 13:25]
  assign io_metadata_init_bits_desc_state_field_type_19_is_host = _T_1 ? 1'h0 : _GEN_1511; // @[Conditional.scala 40:58 Util.scala 13:25]
  assign io_metadata_init_bits_desc_state_field_type_20_is_repeated = _T_1 ? 1'h0 : _GEN_1518; // @[Conditional.scala 40:58 Util.scala 13:25]
  assign io_metadata_init_bits_desc_state_field_type_20_field_type = _T_1 ? 5'h0 : _GEN_1517; // @[Conditional.scala 40:58 Util.scala 13:25]
  assign io_metadata_init_bits_desc_state_field_type_20_sub_class_id = _T_1 ? 16'h0 : _GEN_1516; // @[Conditional.scala 40:58 Util.scala 13:25]
  assign io_metadata_init_bits_desc_state_field_type_20_is_host = _T_1 ? 1'h0 : _GEN_1515; // @[Conditional.scala 40:58 Util.scala 13:25]
  assign io_metadata_init_bits_desc_state_field_type_21_is_repeated = _T_1 ? 1'h0 : _GEN_1522; // @[Conditional.scala 40:58 Util.scala 13:25]
  assign io_metadata_init_bits_desc_state_field_type_21_field_type = _T_1 ? 5'h0 : _GEN_1521; // @[Conditional.scala 40:58 Util.scala 13:25]
  assign io_metadata_init_bits_desc_state_field_type_21_sub_class_id = _T_1 ? 16'h0 : _GEN_1520; // @[Conditional.scala 40:58 Util.scala 13:25]
  assign io_metadata_init_bits_desc_state_field_type_21_is_host = _T_1 ? 1'h0 : _GEN_1519; // @[Conditional.scala 40:58 Util.scala 13:25]
  assign io_metadata_init_bits_desc_state_field_type_22_is_repeated = _T_1 ? 1'h0 : _GEN_1526; // @[Conditional.scala 40:58 Util.scala 13:25]
  assign io_metadata_init_bits_desc_state_field_type_22_field_type = _T_1 ? 5'h0 : _GEN_1525; // @[Conditional.scala 40:58 Util.scala 13:25]
  assign io_metadata_init_bits_desc_state_field_type_22_sub_class_id = _T_1 ? 16'h0 : _GEN_1524; // @[Conditional.scala 40:58 Util.scala 13:25]
  assign io_metadata_init_bits_desc_state_field_type_22_is_host = _T_1 ? 1'h0 : _GEN_1523; // @[Conditional.scala 40:58 Util.scala 13:25]
  assign io_metadata_init_bits_desc_state_field_type_23_is_repeated = _T_1 ? 1'h0 : _GEN_1530; // @[Conditional.scala 40:58 Util.scala 13:25]
  assign io_metadata_init_bits_desc_state_field_type_23_field_type = _T_1 ? 5'h0 : _GEN_1529; // @[Conditional.scala 40:58 Util.scala 13:25]
  assign io_metadata_init_bits_desc_state_field_type_23_sub_class_id = _T_1 ? 16'h0 : _GEN_1528; // @[Conditional.scala 40:58 Util.scala 13:25]
  assign io_metadata_init_bits_desc_state_field_type_23_is_host = _T_1 ? 1'h0 : _GEN_1527; // @[Conditional.scala 40:58 Util.scala 13:25]
  assign io_metadata_init_bits_desc_state_field_type_24_is_repeated = _T_1 ? 1'h0 : _GEN_1534; // @[Conditional.scala 40:58 Util.scala 13:25]
  assign io_metadata_init_bits_desc_state_field_type_24_field_type = _T_1 ? 5'h0 : _GEN_1533; // @[Conditional.scala 40:58 Util.scala 13:25]
  assign io_metadata_init_bits_desc_state_field_type_24_sub_class_id = _T_1 ? 16'h0 : _GEN_1532; // @[Conditional.scala 40:58 Util.scala 13:25]
  assign io_metadata_init_bits_desc_state_field_type_24_is_host = _T_1 ? 1'h0 : _GEN_1531; // @[Conditional.scala 40:58 Util.scala 13:25]
  assign io_metadata_init_bits_desc_state_field_type_25_is_repeated = _T_1 ? 1'h0 : _GEN_1538; // @[Conditional.scala 40:58 Util.scala 13:25]
  assign io_metadata_init_bits_desc_state_field_type_25_field_type = _T_1 ? 5'h0 : _GEN_1537; // @[Conditional.scala 40:58 Util.scala 13:25]
  assign io_metadata_init_bits_desc_state_field_type_25_sub_class_id = _T_1 ? 16'h0 : _GEN_1536; // @[Conditional.scala 40:58 Util.scala 13:25]
  assign io_metadata_init_bits_desc_state_field_type_25_is_host = _T_1 ? 1'h0 : _GEN_1535; // @[Conditional.scala 40:58 Util.scala 13:25]
  assign io_metadata_init_bits_desc_state_field_type_26_is_repeated = _T_1 ? 1'h0 : _GEN_1542; // @[Conditional.scala 40:58 Util.scala 13:25]
  assign io_metadata_init_bits_desc_state_field_type_26_field_type = _T_1 ? 5'h0 : _GEN_1541; // @[Conditional.scala 40:58 Util.scala 13:25]
  assign io_metadata_init_bits_desc_state_field_type_26_sub_class_id = _T_1 ? 16'h0 : _GEN_1540; // @[Conditional.scala 40:58 Util.scala 13:25]
  assign io_metadata_init_bits_desc_state_field_type_26_is_host = _T_1 ? 1'h0 : _GEN_1539; // @[Conditional.scala 40:58 Util.scala 13:25]
  assign io_metadata_init_bits_desc_state_field_type_27_is_repeated = _T_1 ? 1'h0 : _GEN_1546; // @[Conditional.scala 40:58 Util.scala 13:25]
  assign io_metadata_init_bits_desc_state_field_type_27_field_type = _T_1 ? 5'h0 : _GEN_1545; // @[Conditional.scala 40:58 Util.scala 13:25]
  assign io_metadata_init_bits_desc_state_field_type_27_sub_class_id = _T_1 ? 16'h0 : _GEN_1544; // @[Conditional.scala 40:58 Util.scala 13:25]
  assign io_metadata_init_bits_desc_state_field_type_27_is_host = _T_1 ? 1'h0 : _GEN_1543; // @[Conditional.scala 40:58 Util.scala 13:25]
  assign io_metadata_init_bits_desc_state_field_type_28_is_repeated = _T_1 ? 1'h0 : _GEN_1550; // @[Conditional.scala 40:58 Util.scala 13:25]
  assign io_metadata_init_bits_desc_state_field_type_28_field_type = _T_1 ? 5'h0 : _GEN_1549; // @[Conditional.scala 40:58 Util.scala 13:25]
  assign io_metadata_init_bits_desc_state_field_type_28_sub_class_id = _T_1 ? 16'h0 : _GEN_1548; // @[Conditional.scala 40:58 Util.scala 13:25]
  assign io_metadata_init_bits_desc_state_field_type_28_is_host = _T_1 ? 1'h0 : _GEN_1547; // @[Conditional.scala 40:58 Util.scala 13:25]
  assign io_metadata_init_bits_desc_state_field_type_29_is_repeated = _T_1 ? 1'h0 : _GEN_1554; // @[Conditional.scala 40:58 Util.scala 13:25]
  assign io_metadata_init_bits_desc_state_field_type_29_field_type = _T_1 ? 5'h0 : _GEN_1553; // @[Conditional.scala 40:58 Util.scala 13:25]
  assign io_metadata_init_bits_desc_state_field_type_29_sub_class_id = _T_1 ? 16'h0 : _GEN_1552; // @[Conditional.scala 40:58 Util.scala 13:25]
  assign io_metadata_init_bits_desc_state_field_type_29_is_host = _T_1 ? 1'h0 : _GEN_1551; // @[Conditional.scala 40:58 Util.scala 13:25]
  assign io_metadata_init_bits_desc_state_field_type_30_is_repeated = _T_1 ? 1'h0 : _GEN_1558; // @[Conditional.scala 40:58 Util.scala 13:25]
  assign io_metadata_init_bits_desc_state_field_type_30_field_type = _T_1 ? 5'h0 : _GEN_1557; // @[Conditional.scala 40:58 Util.scala 13:25]
  assign io_metadata_init_bits_desc_state_field_type_30_sub_class_id = _T_1 ? 16'h0 : _GEN_1556; // @[Conditional.scala 40:58 Util.scala 13:25]
  assign io_metadata_init_bits_desc_state_field_type_30_is_host = _T_1 ? 1'h0 : _GEN_1555; // @[Conditional.scala 40:58 Util.scala 13:25]
  assign io_metadata_init_bits_desc_state_field_type_31_is_repeated = _T_1 ? 1'h0 : _GEN_1562; // @[Conditional.scala 40:58 Util.scala 13:25]
  assign io_metadata_init_bits_desc_state_field_type_31_field_type = _T_1 ? 5'h0 : _GEN_1561; // @[Conditional.scala 40:58 Util.scala 13:25]
  assign io_metadata_init_bits_desc_state_field_type_31_sub_class_id = _T_1 ? 16'h0 : _GEN_1560; // @[Conditional.scala 40:58 Util.scala 13:25]
  assign io_metadata_init_bits_desc_state_field_type_31_is_host = _T_1 ? 1'h0 : _GEN_1559; // @[Conditional.scala 40:58 Util.scala 13:25]
  assign io_metadata_init_bits_desc_state_field_type_32_is_repeated = _T_1 ? 1'h0 : _GEN_1566; // @[Conditional.scala 40:58 Util.scala 13:25]
  assign io_metadata_init_bits_desc_state_field_type_32_field_type = _T_1 ? 5'h0 : _GEN_1565; // @[Conditional.scala 40:58 Util.scala 13:25]
  assign io_metadata_init_bits_desc_state_field_type_32_sub_class_id = _T_1 ? 16'h0 : _GEN_1564; // @[Conditional.scala 40:58 Util.scala 13:25]
  assign io_metadata_init_bits_desc_state_field_type_32_is_host = _T_1 ? 1'h0 : _GEN_1563; // @[Conditional.scala 40:58 Util.scala 13:25]
  assign io_ser_cmd_valid = _T_1 ? 1'h0 : _GEN_1582; // @[Conditional.scala 40:58 Util.scala 13:25]
  assign io_ser_cmd_bits_class_id = _GEN_1872[9:0];
  assign io_ser_cmd_bits_host_base_addr = _T_1 ? 64'h0 : _GEN_1584; // @[Conditional.scala 40:58 Util.scala 13:25]
  always @(posedge clock) begin
    if (reset) begin // @[Control.scala 43:27]
      s_wr <= 3'h0; // @[Control.scala 43:27]
    end else if (_T_1) begin // @[Conditional.scala 40:58]
      if (_T_2) begin // @[Control.scala 74:40]
        if (_w_addr_T == 64'ha) begin // @[Control.scala 76:84]
          s_wr <= 3'h2; // @[Control.scala 77:33]
        end else begin
          s_wr <= _GEN_5;
        end
      end
    end else if (_T_15) begin // @[Conditional.scala 39:67]
      s_wr <= _GEN_11;
    end else if (_T_17) begin // @[Conditional.scala 39:67]
      s_wr <= _GEN_11;
    end else begin
      s_wr <= _GEN_800;
    end
    if (reset) begin // @[Control.scala 56:31]
      cur_data <= 32'h0; // @[Control.scala 56:31]
    end else if (_T) begin // @[Control.scala 58:23]
      cur_data <= _cur_data_T_1; // @[Control.scala 59:26]
    end
    if (reset) begin // @[Control.scala 57:36]
      classmeta_reg_class_id <= 10'h0; // @[Control.scala 57:36]
    end else begin
      classmeta_reg_class_id <= _GEN_1600[9:0];
    end
    if (reset) begin // @[Control.scala 57:36]
      classmeta_reg_desc_state_class_length <= 16'h0; // @[Control.scala 57:36]
    end else begin
      classmeta_reg_desc_state_class_length <= _GEN_1602[15:0];
    end
    if (reset) begin // @[Control.scala 57:36]
      classmeta_reg_desc_state_max_field_num <= 8'h0; // @[Control.scala 57:36]
    end else begin
      classmeta_reg_desc_state_max_field_num <= _GEN_1601[7:0];
    end
    if (reset) begin // @[Control.scala 57:36]
      classmeta_reg_desc_state_field_type_0_is_repeated <= 1'h0; // @[Control.scala 57:36]
    end else if (!(_T_1)) begin // @[Conditional.scala 40:58]
      if (!(_T_15)) begin // @[Conditional.scala 39:67]
        if (_T_17) begin // @[Conditional.scala 39:67]
          classmeta_reg_desc_state_field_type_0_is_repeated <= _GEN_16;
        end else begin
          classmeta_reg_desc_state_field_type_0_is_repeated <= _GEN_940;
        end
      end
    end
    if (reset) begin // @[Control.scala 57:36]
      classmeta_reg_desc_state_field_type_0_field_type <= 5'h0; // @[Control.scala 57:36]
    end else if (!(_T_1)) begin // @[Conditional.scala 40:58]
      if (!(_T_15)) begin // @[Conditional.scala 39:67]
        if (_T_17) begin // @[Conditional.scala 39:67]
          classmeta_reg_desc_state_field_type_0_field_type <= _GEN_17;
        end else begin
          classmeta_reg_desc_state_field_type_0_field_type <= _GEN_939;
        end
      end
    end
    if (reset) begin // @[Control.scala 57:36]
      classmeta_reg_desc_state_field_type_0_sub_class_id <= 16'h0; // @[Control.scala 57:36]
    end else if (!(_T_1)) begin // @[Conditional.scala 40:58]
      if (!(_T_15)) begin // @[Conditional.scala 39:67]
        if (_T_17) begin // @[Conditional.scala 39:67]
          classmeta_reg_desc_state_field_type_0_sub_class_id <= _GEN_18;
        end else begin
          classmeta_reg_desc_state_field_type_0_sub_class_id <= _GEN_938;
        end
      end
    end
    if (reset) begin // @[Control.scala 57:36]
      classmeta_reg_desc_state_field_type_0_is_host <= 1'h0; // @[Control.scala 57:36]
    end else if (!(_T_1)) begin // @[Conditional.scala 40:58]
      if (!(_T_15)) begin // @[Conditional.scala 39:67]
        if (_T_17) begin // @[Conditional.scala 39:67]
          classmeta_reg_desc_state_field_type_0_is_host <= _GEN_15;
        end else begin
          classmeta_reg_desc_state_field_type_0_is_host <= _GEN_937;
        end
      end
    end
    if (reset) begin // @[Control.scala 57:36]
      classmeta_reg_desc_state_field_type_1_is_repeated <= 1'h0; // @[Control.scala 57:36]
    end else if (!(_T_1)) begin // @[Conditional.scala 40:58]
      if (!(_T_15)) begin // @[Conditional.scala 39:67]
        if (_T_17) begin // @[Conditional.scala 39:67]
          classmeta_reg_desc_state_field_type_1_is_repeated <= _GEN_20;
        end else begin
          classmeta_reg_desc_state_field_type_1_is_repeated <= _GEN_944;
        end
      end
    end
    if (reset) begin // @[Control.scala 57:36]
      classmeta_reg_desc_state_field_type_1_field_type <= 5'h0; // @[Control.scala 57:36]
    end else if (!(_T_1)) begin // @[Conditional.scala 40:58]
      if (!(_T_15)) begin // @[Conditional.scala 39:67]
        if (_T_17) begin // @[Conditional.scala 39:67]
          classmeta_reg_desc_state_field_type_1_field_type <= _GEN_21;
        end else begin
          classmeta_reg_desc_state_field_type_1_field_type <= _GEN_943;
        end
      end
    end
    if (reset) begin // @[Control.scala 57:36]
      classmeta_reg_desc_state_field_type_1_sub_class_id <= 16'h0; // @[Control.scala 57:36]
    end else if (!(_T_1)) begin // @[Conditional.scala 40:58]
      if (!(_T_15)) begin // @[Conditional.scala 39:67]
        if (_T_17) begin // @[Conditional.scala 39:67]
          classmeta_reg_desc_state_field_type_1_sub_class_id <= _GEN_22;
        end else begin
          classmeta_reg_desc_state_field_type_1_sub_class_id <= _GEN_942;
        end
      end
    end
    if (reset) begin // @[Control.scala 57:36]
      classmeta_reg_desc_state_field_type_1_is_host <= 1'h0; // @[Control.scala 57:36]
    end else if (!(_T_1)) begin // @[Conditional.scala 40:58]
      if (!(_T_15)) begin // @[Conditional.scala 39:67]
        if (_T_17) begin // @[Conditional.scala 39:67]
          classmeta_reg_desc_state_field_type_1_is_host <= _GEN_19;
        end else begin
          classmeta_reg_desc_state_field_type_1_is_host <= _GEN_941;
        end
      end
    end
    if (reset) begin // @[Control.scala 57:36]
      classmeta_reg_desc_state_field_type_2_is_repeated <= 1'h0; // @[Control.scala 57:36]
    end else if (!(_T_1)) begin // @[Conditional.scala 40:58]
      if (!(_T_15)) begin // @[Conditional.scala 39:67]
        if (_T_17) begin // @[Conditional.scala 39:67]
          classmeta_reg_desc_state_field_type_2_is_repeated <= _GEN_24;
        end else begin
          classmeta_reg_desc_state_field_type_2_is_repeated <= _GEN_948;
        end
      end
    end
    if (reset) begin // @[Control.scala 57:36]
      classmeta_reg_desc_state_field_type_2_field_type <= 5'h0; // @[Control.scala 57:36]
    end else if (!(_T_1)) begin // @[Conditional.scala 40:58]
      if (!(_T_15)) begin // @[Conditional.scala 39:67]
        if (_T_17) begin // @[Conditional.scala 39:67]
          classmeta_reg_desc_state_field_type_2_field_type <= _GEN_25;
        end else begin
          classmeta_reg_desc_state_field_type_2_field_type <= _GEN_947;
        end
      end
    end
    if (reset) begin // @[Control.scala 57:36]
      classmeta_reg_desc_state_field_type_2_sub_class_id <= 16'h0; // @[Control.scala 57:36]
    end else if (!(_T_1)) begin // @[Conditional.scala 40:58]
      if (!(_T_15)) begin // @[Conditional.scala 39:67]
        if (_T_17) begin // @[Conditional.scala 39:67]
          classmeta_reg_desc_state_field_type_2_sub_class_id <= _GEN_26;
        end else begin
          classmeta_reg_desc_state_field_type_2_sub_class_id <= _GEN_946;
        end
      end
    end
    if (reset) begin // @[Control.scala 57:36]
      classmeta_reg_desc_state_field_type_2_is_host <= 1'h0; // @[Control.scala 57:36]
    end else if (!(_T_1)) begin // @[Conditional.scala 40:58]
      if (!(_T_15)) begin // @[Conditional.scala 39:67]
        if (_T_17) begin // @[Conditional.scala 39:67]
          classmeta_reg_desc_state_field_type_2_is_host <= _GEN_23;
        end else begin
          classmeta_reg_desc_state_field_type_2_is_host <= _GEN_945;
        end
      end
    end
    if (reset) begin // @[Control.scala 57:36]
      classmeta_reg_desc_state_field_type_3_is_repeated <= 1'h0; // @[Control.scala 57:36]
    end else if (!(_T_1)) begin // @[Conditional.scala 40:58]
      if (!(_T_15)) begin // @[Conditional.scala 39:67]
        if (_T_17) begin // @[Conditional.scala 39:67]
          classmeta_reg_desc_state_field_type_3_is_repeated <= _GEN_28;
        end else begin
          classmeta_reg_desc_state_field_type_3_is_repeated <= _GEN_952;
        end
      end
    end
    if (reset) begin // @[Control.scala 57:36]
      classmeta_reg_desc_state_field_type_3_field_type <= 5'h0; // @[Control.scala 57:36]
    end else if (!(_T_1)) begin // @[Conditional.scala 40:58]
      if (!(_T_15)) begin // @[Conditional.scala 39:67]
        if (_T_17) begin // @[Conditional.scala 39:67]
          classmeta_reg_desc_state_field_type_3_field_type <= _GEN_29;
        end else begin
          classmeta_reg_desc_state_field_type_3_field_type <= _GEN_951;
        end
      end
    end
    if (reset) begin // @[Control.scala 57:36]
      classmeta_reg_desc_state_field_type_3_sub_class_id <= 16'h0; // @[Control.scala 57:36]
    end else if (!(_T_1)) begin // @[Conditional.scala 40:58]
      if (!(_T_15)) begin // @[Conditional.scala 39:67]
        if (_T_17) begin // @[Conditional.scala 39:67]
          classmeta_reg_desc_state_field_type_3_sub_class_id <= _GEN_30;
        end else begin
          classmeta_reg_desc_state_field_type_3_sub_class_id <= _GEN_950;
        end
      end
    end
    if (reset) begin // @[Control.scala 57:36]
      classmeta_reg_desc_state_field_type_3_is_host <= 1'h0; // @[Control.scala 57:36]
    end else if (!(_T_1)) begin // @[Conditional.scala 40:58]
      if (!(_T_15)) begin // @[Conditional.scala 39:67]
        if (_T_17) begin // @[Conditional.scala 39:67]
          classmeta_reg_desc_state_field_type_3_is_host <= _GEN_27;
        end else begin
          classmeta_reg_desc_state_field_type_3_is_host <= _GEN_949;
        end
      end
    end
    if (reset) begin // @[Control.scala 57:36]
      classmeta_reg_desc_state_field_type_4_is_repeated <= 1'h0; // @[Control.scala 57:36]
    end else if (!(_T_1)) begin // @[Conditional.scala 40:58]
      if (!(_T_15)) begin // @[Conditional.scala 39:67]
        if (_T_17) begin // @[Conditional.scala 39:67]
          classmeta_reg_desc_state_field_type_4_is_repeated <= _GEN_32;
        end else begin
          classmeta_reg_desc_state_field_type_4_is_repeated <= _GEN_956;
        end
      end
    end
    if (reset) begin // @[Control.scala 57:36]
      classmeta_reg_desc_state_field_type_4_field_type <= 5'h0; // @[Control.scala 57:36]
    end else if (!(_T_1)) begin // @[Conditional.scala 40:58]
      if (!(_T_15)) begin // @[Conditional.scala 39:67]
        if (_T_17) begin // @[Conditional.scala 39:67]
          classmeta_reg_desc_state_field_type_4_field_type <= _GEN_33;
        end else begin
          classmeta_reg_desc_state_field_type_4_field_type <= _GEN_955;
        end
      end
    end
    if (reset) begin // @[Control.scala 57:36]
      classmeta_reg_desc_state_field_type_4_sub_class_id <= 16'h0; // @[Control.scala 57:36]
    end else if (!(_T_1)) begin // @[Conditional.scala 40:58]
      if (!(_T_15)) begin // @[Conditional.scala 39:67]
        if (_T_17) begin // @[Conditional.scala 39:67]
          classmeta_reg_desc_state_field_type_4_sub_class_id <= _GEN_34;
        end else begin
          classmeta_reg_desc_state_field_type_4_sub_class_id <= _GEN_954;
        end
      end
    end
    if (reset) begin // @[Control.scala 57:36]
      classmeta_reg_desc_state_field_type_4_is_host <= 1'h0; // @[Control.scala 57:36]
    end else if (!(_T_1)) begin // @[Conditional.scala 40:58]
      if (!(_T_15)) begin // @[Conditional.scala 39:67]
        if (_T_17) begin // @[Conditional.scala 39:67]
          classmeta_reg_desc_state_field_type_4_is_host <= _GEN_31;
        end else begin
          classmeta_reg_desc_state_field_type_4_is_host <= _GEN_953;
        end
      end
    end
    if (reset) begin // @[Control.scala 57:36]
      classmeta_reg_desc_state_field_type_5_is_repeated <= 1'h0; // @[Control.scala 57:36]
    end else if (!(_T_1)) begin // @[Conditional.scala 40:58]
      if (!(_T_15)) begin // @[Conditional.scala 39:67]
        if (_T_17) begin // @[Conditional.scala 39:67]
          classmeta_reg_desc_state_field_type_5_is_repeated <= _GEN_36;
        end else begin
          classmeta_reg_desc_state_field_type_5_is_repeated <= _GEN_960;
        end
      end
    end
    if (reset) begin // @[Control.scala 57:36]
      classmeta_reg_desc_state_field_type_5_field_type <= 5'h0; // @[Control.scala 57:36]
    end else if (!(_T_1)) begin // @[Conditional.scala 40:58]
      if (!(_T_15)) begin // @[Conditional.scala 39:67]
        if (_T_17) begin // @[Conditional.scala 39:67]
          classmeta_reg_desc_state_field_type_5_field_type <= _GEN_37;
        end else begin
          classmeta_reg_desc_state_field_type_5_field_type <= _GEN_959;
        end
      end
    end
    if (reset) begin // @[Control.scala 57:36]
      classmeta_reg_desc_state_field_type_5_sub_class_id <= 16'h0; // @[Control.scala 57:36]
    end else if (!(_T_1)) begin // @[Conditional.scala 40:58]
      if (!(_T_15)) begin // @[Conditional.scala 39:67]
        if (_T_17) begin // @[Conditional.scala 39:67]
          classmeta_reg_desc_state_field_type_5_sub_class_id <= _GEN_38;
        end else begin
          classmeta_reg_desc_state_field_type_5_sub_class_id <= _GEN_958;
        end
      end
    end
    if (reset) begin // @[Control.scala 57:36]
      classmeta_reg_desc_state_field_type_5_is_host <= 1'h0; // @[Control.scala 57:36]
    end else if (!(_T_1)) begin // @[Conditional.scala 40:58]
      if (!(_T_15)) begin // @[Conditional.scala 39:67]
        if (_T_17) begin // @[Conditional.scala 39:67]
          classmeta_reg_desc_state_field_type_5_is_host <= _GEN_35;
        end else begin
          classmeta_reg_desc_state_field_type_5_is_host <= _GEN_957;
        end
      end
    end
    if (reset) begin // @[Control.scala 57:36]
      classmeta_reg_desc_state_field_type_6_is_repeated <= 1'h0; // @[Control.scala 57:36]
    end else if (!(_T_1)) begin // @[Conditional.scala 40:58]
      if (!(_T_15)) begin // @[Conditional.scala 39:67]
        if (_T_17) begin // @[Conditional.scala 39:67]
          classmeta_reg_desc_state_field_type_6_is_repeated <= _GEN_40;
        end else begin
          classmeta_reg_desc_state_field_type_6_is_repeated <= _GEN_964;
        end
      end
    end
    if (reset) begin // @[Control.scala 57:36]
      classmeta_reg_desc_state_field_type_6_field_type <= 5'h0; // @[Control.scala 57:36]
    end else if (!(_T_1)) begin // @[Conditional.scala 40:58]
      if (!(_T_15)) begin // @[Conditional.scala 39:67]
        if (_T_17) begin // @[Conditional.scala 39:67]
          classmeta_reg_desc_state_field_type_6_field_type <= _GEN_41;
        end else begin
          classmeta_reg_desc_state_field_type_6_field_type <= _GEN_963;
        end
      end
    end
    if (reset) begin // @[Control.scala 57:36]
      classmeta_reg_desc_state_field_type_6_sub_class_id <= 16'h0; // @[Control.scala 57:36]
    end else if (!(_T_1)) begin // @[Conditional.scala 40:58]
      if (!(_T_15)) begin // @[Conditional.scala 39:67]
        if (_T_17) begin // @[Conditional.scala 39:67]
          classmeta_reg_desc_state_field_type_6_sub_class_id <= _GEN_42;
        end else begin
          classmeta_reg_desc_state_field_type_6_sub_class_id <= _GEN_962;
        end
      end
    end
    if (reset) begin // @[Control.scala 57:36]
      classmeta_reg_desc_state_field_type_6_is_host <= 1'h0; // @[Control.scala 57:36]
    end else if (!(_T_1)) begin // @[Conditional.scala 40:58]
      if (!(_T_15)) begin // @[Conditional.scala 39:67]
        if (_T_17) begin // @[Conditional.scala 39:67]
          classmeta_reg_desc_state_field_type_6_is_host <= _GEN_39;
        end else begin
          classmeta_reg_desc_state_field_type_6_is_host <= _GEN_961;
        end
      end
    end
    if (reset) begin // @[Control.scala 57:36]
      classmeta_reg_desc_state_field_type_7_is_repeated <= 1'h0; // @[Control.scala 57:36]
    end else if (!(_T_1)) begin // @[Conditional.scala 40:58]
      if (!(_T_15)) begin // @[Conditional.scala 39:67]
        if (_T_17) begin // @[Conditional.scala 39:67]
          classmeta_reg_desc_state_field_type_7_is_repeated <= _GEN_44;
        end else begin
          classmeta_reg_desc_state_field_type_7_is_repeated <= _GEN_968;
        end
      end
    end
    if (reset) begin // @[Control.scala 57:36]
      classmeta_reg_desc_state_field_type_7_field_type <= 5'h0; // @[Control.scala 57:36]
    end else if (!(_T_1)) begin // @[Conditional.scala 40:58]
      if (!(_T_15)) begin // @[Conditional.scala 39:67]
        if (_T_17) begin // @[Conditional.scala 39:67]
          classmeta_reg_desc_state_field_type_7_field_type <= _GEN_45;
        end else begin
          classmeta_reg_desc_state_field_type_7_field_type <= _GEN_967;
        end
      end
    end
    if (reset) begin // @[Control.scala 57:36]
      classmeta_reg_desc_state_field_type_7_sub_class_id <= 16'h0; // @[Control.scala 57:36]
    end else if (!(_T_1)) begin // @[Conditional.scala 40:58]
      if (!(_T_15)) begin // @[Conditional.scala 39:67]
        if (_T_17) begin // @[Conditional.scala 39:67]
          classmeta_reg_desc_state_field_type_7_sub_class_id <= _GEN_46;
        end else begin
          classmeta_reg_desc_state_field_type_7_sub_class_id <= _GEN_966;
        end
      end
    end
    if (reset) begin // @[Control.scala 57:36]
      classmeta_reg_desc_state_field_type_7_is_host <= 1'h0; // @[Control.scala 57:36]
    end else if (!(_T_1)) begin // @[Conditional.scala 40:58]
      if (!(_T_15)) begin // @[Conditional.scala 39:67]
        if (_T_17) begin // @[Conditional.scala 39:67]
          classmeta_reg_desc_state_field_type_7_is_host <= _GEN_43;
        end else begin
          classmeta_reg_desc_state_field_type_7_is_host <= _GEN_965;
        end
      end
    end
    if (reset) begin // @[Control.scala 57:36]
      classmeta_reg_desc_state_field_type_8_is_repeated <= 1'h0; // @[Control.scala 57:36]
    end else if (!(_T_1)) begin // @[Conditional.scala 40:58]
      if (!(_T_15)) begin // @[Conditional.scala 39:67]
        if (_T_17) begin // @[Conditional.scala 39:67]
          classmeta_reg_desc_state_field_type_8_is_repeated <= _GEN_48;
        end else begin
          classmeta_reg_desc_state_field_type_8_is_repeated <= _GEN_972;
        end
      end
    end
    if (reset) begin // @[Control.scala 57:36]
      classmeta_reg_desc_state_field_type_8_field_type <= 5'h0; // @[Control.scala 57:36]
    end else if (!(_T_1)) begin // @[Conditional.scala 40:58]
      if (!(_T_15)) begin // @[Conditional.scala 39:67]
        if (_T_17) begin // @[Conditional.scala 39:67]
          classmeta_reg_desc_state_field_type_8_field_type <= _GEN_49;
        end else begin
          classmeta_reg_desc_state_field_type_8_field_type <= _GEN_971;
        end
      end
    end
    if (reset) begin // @[Control.scala 57:36]
      classmeta_reg_desc_state_field_type_8_sub_class_id <= 16'h0; // @[Control.scala 57:36]
    end else if (!(_T_1)) begin // @[Conditional.scala 40:58]
      if (!(_T_15)) begin // @[Conditional.scala 39:67]
        if (_T_17) begin // @[Conditional.scala 39:67]
          classmeta_reg_desc_state_field_type_8_sub_class_id <= _GEN_50;
        end else begin
          classmeta_reg_desc_state_field_type_8_sub_class_id <= _GEN_970;
        end
      end
    end
    if (reset) begin // @[Control.scala 57:36]
      classmeta_reg_desc_state_field_type_8_is_host <= 1'h0; // @[Control.scala 57:36]
    end else if (!(_T_1)) begin // @[Conditional.scala 40:58]
      if (!(_T_15)) begin // @[Conditional.scala 39:67]
        if (_T_17) begin // @[Conditional.scala 39:67]
          classmeta_reg_desc_state_field_type_8_is_host <= _GEN_47;
        end else begin
          classmeta_reg_desc_state_field_type_8_is_host <= _GEN_969;
        end
      end
    end
    if (reset) begin // @[Control.scala 57:36]
      classmeta_reg_desc_state_field_type_9_is_repeated <= 1'h0; // @[Control.scala 57:36]
    end else if (!(_T_1)) begin // @[Conditional.scala 40:58]
      if (!(_T_15)) begin // @[Conditional.scala 39:67]
        if (_T_17) begin // @[Conditional.scala 39:67]
          classmeta_reg_desc_state_field_type_9_is_repeated <= _GEN_52;
        end else begin
          classmeta_reg_desc_state_field_type_9_is_repeated <= _GEN_976;
        end
      end
    end
    if (reset) begin // @[Control.scala 57:36]
      classmeta_reg_desc_state_field_type_9_field_type <= 5'h0; // @[Control.scala 57:36]
    end else if (!(_T_1)) begin // @[Conditional.scala 40:58]
      if (!(_T_15)) begin // @[Conditional.scala 39:67]
        if (_T_17) begin // @[Conditional.scala 39:67]
          classmeta_reg_desc_state_field_type_9_field_type <= _GEN_53;
        end else begin
          classmeta_reg_desc_state_field_type_9_field_type <= _GEN_975;
        end
      end
    end
    if (reset) begin // @[Control.scala 57:36]
      classmeta_reg_desc_state_field_type_9_sub_class_id <= 16'h0; // @[Control.scala 57:36]
    end else if (!(_T_1)) begin // @[Conditional.scala 40:58]
      if (!(_T_15)) begin // @[Conditional.scala 39:67]
        if (_T_17) begin // @[Conditional.scala 39:67]
          classmeta_reg_desc_state_field_type_9_sub_class_id <= _GEN_54;
        end else begin
          classmeta_reg_desc_state_field_type_9_sub_class_id <= _GEN_974;
        end
      end
    end
    if (reset) begin // @[Control.scala 57:36]
      classmeta_reg_desc_state_field_type_9_is_host <= 1'h0; // @[Control.scala 57:36]
    end else if (!(_T_1)) begin // @[Conditional.scala 40:58]
      if (!(_T_15)) begin // @[Conditional.scala 39:67]
        if (_T_17) begin // @[Conditional.scala 39:67]
          classmeta_reg_desc_state_field_type_9_is_host <= _GEN_51;
        end else begin
          classmeta_reg_desc_state_field_type_9_is_host <= _GEN_973;
        end
      end
    end
    if (reset) begin // @[Control.scala 57:36]
      classmeta_reg_desc_state_field_type_10_is_repeated <= 1'h0; // @[Control.scala 57:36]
    end else if (!(_T_1)) begin // @[Conditional.scala 40:58]
      if (!(_T_15)) begin // @[Conditional.scala 39:67]
        if (_T_17) begin // @[Conditional.scala 39:67]
          classmeta_reg_desc_state_field_type_10_is_repeated <= _GEN_56;
        end else begin
          classmeta_reg_desc_state_field_type_10_is_repeated <= _GEN_980;
        end
      end
    end
    if (reset) begin // @[Control.scala 57:36]
      classmeta_reg_desc_state_field_type_10_field_type <= 5'h0; // @[Control.scala 57:36]
    end else if (!(_T_1)) begin // @[Conditional.scala 40:58]
      if (!(_T_15)) begin // @[Conditional.scala 39:67]
        if (_T_17) begin // @[Conditional.scala 39:67]
          classmeta_reg_desc_state_field_type_10_field_type <= _GEN_57;
        end else begin
          classmeta_reg_desc_state_field_type_10_field_type <= _GEN_979;
        end
      end
    end
    if (reset) begin // @[Control.scala 57:36]
      classmeta_reg_desc_state_field_type_10_sub_class_id <= 16'h0; // @[Control.scala 57:36]
    end else if (!(_T_1)) begin // @[Conditional.scala 40:58]
      if (!(_T_15)) begin // @[Conditional.scala 39:67]
        if (_T_17) begin // @[Conditional.scala 39:67]
          classmeta_reg_desc_state_field_type_10_sub_class_id <= _GEN_58;
        end else begin
          classmeta_reg_desc_state_field_type_10_sub_class_id <= _GEN_978;
        end
      end
    end
    if (reset) begin // @[Control.scala 57:36]
      classmeta_reg_desc_state_field_type_10_is_host <= 1'h0; // @[Control.scala 57:36]
    end else if (!(_T_1)) begin // @[Conditional.scala 40:58]
      if (!(_T_15)) begin // @[Conditional.scala 39:67]
        if (_T_17) begin // @[Conditional.scala 39:67]
          classmeta_reg_desc_state_field_type_10_is_host <= _GEN_55;
        end else begin
          classmeta_reg_desc_state_field_type_10_is_host <= _GEN_977;
        end
      end
    end
    if (reset) begin // @[Control.scala 57:36]
      classmeta_reg_desc_state_field_type_11_is_repeated <= 1'h0; // @[Control.scala 57:36]
    end else if (!(_T_1)) begin // @[Conditional.scala 40:58]
      if (!(_T_15)) begin // @[Conditional.scala 39:67]
        if (_T_17) begin // @[Conditional.scala 39:67]
          classmeta_reg_desc_state_field_type_11_is_repeated <= _GEN_60;
        end else begin
          classmeta_reg_desc_state_field_type_11_is_repeated <= _GEN_984;
        end
      end
    end
    if (reset) begin // @[Control.scala 57:36]
      classmeta_reg_desc_state_field_type_11_field_type <= 5'h0; // @[Control.scala 57:36]
    end else if (!(_T_1)) begin // @[Conditional.scala 40:58]
      if (!(_T_15)) begin // @[Conditional.scala 39:67]
        if (_T_17) begin // @[Conditional.scala 39:67]
          classmeta_reg_desc_state_field_type_11_field_type <= _GEN_61;
        end else begin
          classmeta_reg_desc_state_field_type_11_field_type <= _GEN_983;
        end
      end
    end
    if (reset) begin // @[Control.scala 57:36]
      classmeta_reg_desc_state_field_type_11_sub_class_id <= 16'h0; // @[Control.scala 57:36]
    end else if (!(_T_1)) begin // @[Conditional.scala 40:58]
      if (!(_T_15)) begin // @[Conditional.scala 39:67]
        if (_T_17) begin // @[Conditional.scala 39:67]
          classmeta_reg_desc_state_field_type_11_sub_class_id <= _GEN_62;
        end else begin
          classmeta_reg_desc_state_field_type_11_sub_class_id <= _GEN_982;
        end
      end
    end
    if (reset) begin // @[Control.scala 57:36]
      classmeta_reg_desc_state_field_type_11_is_host <= 1'h0; // @[Control.scala 57:36]
    end else if (!(_T_1)) begin // @[Conditional.scala 40:58]
      if (!(_T_15)) begin // @[Conditional.scala 39:67]
        if (_T_17) begin // @[Conditional.scala 39:67]
          classmeta_reg_desc_state_field_type_11_is_host <= _GEN_59;
        end else begin
          classmeta_reg_desc_state_field_type_11_is_host <= _GEN_981;
        end
      end
    end
    if (reset) begin // @[Control.scala 57:36]
      classmeta_reg_desc_state_field_type_12_is_repeated <= 1'h0; // @[Control.scala 57:36]
    end else if (!(_T_1)) begin // @[Conditional.scala 40:58]
      if (!(_T_15)) begin // @[Conditional.scala 39:67]
        if (_T_17) begin // @[Conditional.scala 39:67]
          classmeta_reg_desc_state_field_type_12_is_repeated <= _GEN_64;
        end else begin
          classmeta_reg_desc_state_field_type_12_is_repeated <= _GEN_988;
        end
      end
    end
    if (reset) begin // @[Control.scala 57:36]
      classmeta_reg_desc_state_field_type_12_field_type <= 5'h0; // @[Control.scala 57:36]
    end else if (!(_T_1)) begin // @[Conditional.scala 40:58]
      if (!(_T_15)) begin // @[Conditional.scala 39:67]
        if (_T_17) begin // @[Conditional.scala 39:67]
          classmeta_reg_desc_state_field_type_12_field_type <= _GEN_65;
        end else begin
          classmeta_reg_desc_state_field_type_12_field_type <= _GEN_987;
        end
      end
    end
    if (reset) begin // @[Control.scala 57:36]
      classmeta_reg_desc_state_field_type_12_sub_class_id <= 16'h0; // @[Control.scala 57:36]
    end else if (!(_T_1)) begin // @[Conditional.scala 40:58]
      if (!(_T_15)) begin // @[Conditional.scala 39:67]
        if (_T_17) begin // @[Conditional.scala 39:67]
          classmeta_reg_desc_state_field_type_12_sub_class_id <= _GEN_66;
        end else begin
          classmeta_reg_desc_state_field_type_12_sub_class_id <= _GEN_986;
        end
      end
    end
    if (reset) begin // @[Control.scala 57:36]
      classmeta_reg_desc_state_field_type_12_is_host <= 1'h0; // @[Control.scala 57:36]
    end else if (!(_T_1)) begin // @[Conditional.scala 40:58]
      if (!(_T_15)) begin // @[Conditional.scala 39:67]
        if (_T_17) begin // @[Conditional.scala 39:67]
          classmeta_reg_desc_state_field_type_12_is_host <= _GEN_63;
        end else begin
          classmeta_reg_desc_state_field_type_12_is_host <= _GEN_985;
        end
      end
    end
    if (reset) begin // @[Control.scala 57:36]
      classmeta_reg_desc_state_field_type_13_is_repeated <= 1'h0; // @[Control.scala 57:36]
    end else if (!(_T_1)) begin // @[Conditional.scala 40:58]
      if (!(_T_15)) begin // @[Conditional.scala 39:67]
        if (_T_17) begin // @[Conditional.scala 39:67]
          classmeta_reg_desc_state_field_type_13_is_repeated <= _GEN_68;
        end else begin
          classmeta_reg_desc_state_field_type_13_is_repeated <= _GEN_992;
        end
      end
    end
    if (reset) begin // @[Control.scala 57:36]
      classmeta_reg_desc_state_field_type_13_field_type <= 5'h0; // @[Control.scala 57:36]
    end else if (!(_T_1)) begin // @[Conditional.scala 40:58]
      if (!(_T_15)) begin // @[Conditional.scala 39:67]
        if (_T_17) begin // @[Conditional.scala 39:67]
          classmeta_reg_desc_state_field_type_13_field_type <= _GEN_69;
        end else begin
          classmeta_reg_desc_state_field_type_13_field_type <= _GEN_991;
        end
      end
    end
    if (reset) begin // @[Control.scala 57:36]
      classmeta_reg_desc_state_field_type_13_sub_class_id <= 16'h0; // @[Control.scala 57:36]
    end else if (!(_T_1)) begin // @[Conditional.scala 40:58]
      if (!(_T_15)) begin // @[Conditional.scala 39:67]
        if (_T_17) begin // @[Conditional.scala 39:67]
          classmeta_reg_desc_state_field_type_13_sub_class_id <= _GEN_70;
        end else begin
          classmeta_reg_desc_state_field_type_13_sub_class_id <= _GEN_990;
        end
      end
    end
    if (reset) begin // @[Control.scala 57:36]
      classmeta_reg_desc_state_field_type_13_is_host <= 1'h0; // @[Control.scala 57:36]
    end else if (!(_T_1)) begin // @[Conditional.scala 40:58]
      if (!(_T_15)) begin // @[Conditional.scala 39:67]
        if (_T_17) begin // @[Conditional.scala 39:67]
          classmeta_reg_desc_state_field_type_13_is_host <= _GEN_67;
        end else begin
          classmeta_reg_desc_state_field_type_13_is_host <= _GEN_989;
        end
      end
    end
    if (reset) begin // @[Control.scala 57:36]
      classmeta_reg_desc_state_field_type_14_is_repeated <= 1'h0; // @[Control.scala 57:36]
    end else if (!(_T_1)) begin // @[Conditional.scala 40:58]
      if (!(_T_15)) begin // @[Conditional.scala 39:67]
        if (!(_T_17)) begin // @[Conditional.scala 39:67]
          classmeta_reg_desc_state_field_type_14_is_repeated <= _GEN_737;
        end
      end
    end
    if (reset) begin // @[Control.scala 57:36]
      classmeta_reg_desc_state_field_type_14_field_type <= 5'h0; // @[Control.scala 57:36]
    end else if (!(_T_1)) begin // @[Conditional.scala 40:58]
      if (!(_T_15)) begin // @[Conditional.scala 39:67]
        if (!(_T_17)) begin // @[Conditional.scala 39:67]
          classmeta_reg_desc_state_field_type_14_field_type <= _GEN_738;
        end
      end
    end
    if (reset) begin // @[Control.scala 57:36]
      classmeta_reg_desc_state_field_type_14_sub_class_id <= 16'h0; // @[Control.scala 57:36]
    end else if (!(_T_1)) begin // @[Conditional.scala 40:58]
      if (!(_T_15)) begin // @[Conditional.scala 39:67]
        if (!(_T_17)) begin // @[Conditional.scala 39:67]
          classmeta_reg_desc_state_field_type_14_sub_class_id <= _GEN_739;
        end
      end
    end
    if (reset) begin // @[Control.scala 57:36]
      classmeta_reg_desc_state_field_type_14_is_host <= 1'h0; // @[Control.scala 57:36]
    end else if (!(_T_1)) begin // @[Conditional.scala 40:58]
      if (!(_T_15)) begin // @[Conditional.scala 39:67]
        if (!(_T_17)) begin // @[Conditional.scala 39:67]
          classmeta_reg_desc_state_field_type_14_is_host <= _GEN_736;
        end
      end
    end
    if (reset) begin // @[Control.scala 57:36]
      classmeta_reg_desc_state_field_type_15_is_repeated <= 1'h0; // @[Control.scala 57:36]
    end else if (!(_T_1)) begin // @[Conditional.scala 40:58]
      if (!(_T_15)) begin // @[Conditional.scala 39:67]
        if (!(_T_17)) begin // @[Conditional.scala 39:67]
          classmeta_reg_desc_state_field_type_15_is_repeated <= _GEN_741;
        end
      end
    end
    if (reset) begin // @[Control.scala 57:36]
      classmeta_reg_desc_state_field_type_15_field_type <= 5'h0; // @[Control.scala 57:36]
    end else if (!(_T_1)) begin // @[Conditional.scala 40:58]
      if (!(_T_15)) begin // @[Conditional.scala 39:67]
        if (!(_T_17)) begin // @[Conditional.scala 39:67]
          classmeta_reg_desc_state_field_type_15_field_type <= _GEN_742;
        end
      end
    end
    if (reset) begin // @[Control.scala 57:36]
      classmeta_reg_desc_state_field_type_15_sub_class_id <= 16'h0; // @[Control.scala 57:36]
    end else if (!(_T_1)) begin // @[Conditional.scala 40:58]
      if (!(_T_15)) begin // @[Conditional.scala 39:67]
        if (!(_T_17)) begin // @[Conditional.scala 39:67]
          classmeta_reg_desc_state_field_type_15_sub_class_id <= _GEN_743;
        end
      end
    end
    if (reset) begin // @[Control.scala 57:36]
      classmeta_reg_desc_state_field_type_15_is_host <= 1'h0; // @[Control.scala 57:36]
    end else if (!(_T_1)) begin // @[Conditional.scala 40:58]
      if (!(_T_15)) begin // @[Conditional.scala 39:67]
        if (!(_T_17)) begin // @[Conditional.scala 39:67]
          classmeta_reg_desc_state_field_type_15_is_host <= _GEN_740;
        end
      end
    end
    if (reset) begin // @[Control.scala 57:36]
      classmeta_reg_desc_state_field_type_16_is_repeated <= 1'h0; // @[Control.scala 57:36]
    end else if (!(_T_1)) begin // @[Conditional.scala 40:58]
      if (!(_T_15)) begin // @[Conditional.scala 39:67]
        if (!(_T_17)) begin // @[Conditional.scala 39:67]
          classmeta_reg_desc_state_field_type_16_is_repeated <= _GEN_745;
        end
      end
    end
    if (reset) begin // @[Control.scala 57:36]
      classmeta_reg_desc_state_field_type_16_field_type <= 5'h0; // @[Control.scala 57:36]
    end else if (!(_T_1)) begin // @[Conditional.scala 40:58]
      if (!(_T_15)) begin // @[Conditional.scala 39:67]
        if (!(_T_17)) begin // @[Conditional.scala 39:67]
          classmeta_reg_desc_state_field_type_16_field_type <= _GEN_746;
        end
      end
    end
    if (reset) begin // @[Control.scala 57:36]
      classmeta_reg_desc_state_field_type_16_sub_class_id <= 16'h0; // @[Control.scala 57:36]
    end else if (!(_T_1)) begin // @[Conditional.scala 40:58]
      if (!(_T_15)) begin // @[Conditional.scala 39:67]
        if (!(_T_17)) begin // @[Conditional.scala 39:67]
          classmeta_reg_desc_state_field_type_16_sub_class_id <= _GEN_747;
        end
      end
    end
    if (reset) begin // @[Control.scala 57:36]
      classmeta_reg_desc_state_field_type_16_is_host <= 1'h0; // @[Control.scala 57:36]
    end else if (!(_T_1)) begin // @[Conditional.scala 40:58]
      if (!(_T_15)) begin // @[Conditional.scala 39:67]
        if (!(_T_17)) begin // @[Conditional.scala 39:67]
          classmeta_reg_desc_state_field_type_16_is_host <= _GEN_744;
        end
      end
    end
    if (reset) begin // @[Control.scala 57:36]
      classmeta_reg_desc_state_field_type_17_is_repeated <= 1'h0; // @[Control.scala 57:36]
    end else if (!(_T_1)) begin // @[Conditional.scala 40:58]
      if (!(_T_15)) begin // @[Conditional.scala 39:67]
        if (!(_T_17)) begin // @[Conditional.scala 39:67]
          classmeta_reg_desc_state_field_type_17_is_repeated <= _GEN_749;
        end
      end
    end
    if (reset) begin // @[Control.scala 57:36]
      classmeta_reg_desc_state_field_type_17_field_type <= 5'h0; // @[Control.scala 57:36]
    end else if (!(_T_1)) begin // @[Conditional.scala 40:58]
      if (!(_T_15)) begin // @[Conditional.scala 39:67]
        if (!(_T_17)) begin // @[Conditional.scala 39:67]
          classmeta_reg_desc_state_field_type_17_field_type <= _GEN_750;
        end
      end
    end
    if (reset) begin // @[Control.scala 57:36]
      classmeta_reg_desc_state_field_type_17_sub_class_id <= 16'h0; // @[Control.scala 57:36]
    end else if (!(_T_1)) begin // @[Conditional.scala 40:58]
      if (!(_T_15)) begin // @[Conditional.scala 39:67]
        if (!(_T_17)) begin // @[Conditional.scala 39:67]
          classmeta_reg_desc_state_field_type_17_sub_class_id <= _GEN_751;
        end
      end
    end
    if (reset) begin // @[Control.scala 57:36]
      classmeta_reg_desc_state_field_type_17_is_host <= 1'h0; // @[Control.scala 57:36]
    end else if (!(_T_1)) begin // @[Conditional.scala 40:58]
      if (!(_T_15)) begin // @[Conditional.scala 39:67]
        if (!(_T_17)) begin // @[Conditional.scala 39:67]
          classmeta_reg_desc_state_field_type_17_is_host <= _GEN_748;
        end
      end
    end
    if (reset) begin // @[Control.scala 57:36]
      classmeta_reg_desc_state_field_type_18_is_repeated <= 1'h0; // @[Control.scala 57:36]
    end else if (!(_T_1)) begin // @[Conditional.scala 40:58]
      if (!(_T_15)) begin // @[Conditional.scala 39:67]
        if (!(_T_17)) begin // @[Conditional.scala 39:67]
          classmeta_reg_desc_state_field_type_18_is_repeated <= _GEN_753;
        end
      end
    end
    if (reset) begin // @[Control.scala 57:36]
      classmeta_reg_desc_state_field_type_18_field_type <= 5'h0; // @[Control.scala 57:36]
    end else if (!(_T_1)) begin // @[Conditional.scala 40:58]
      if (!(_T_15)) begin // @[Conditional.scala 39:67]
        if (!(_T_17)) begin // @[Conditional.scala 39:67]
          classmeta_reg_desc_state_field_type_18_field_type <= _GEN_754;
        end
      end
    end
    if (reset) begin // @[Control.scala 57:36]
      classmeta_reg_desc_state_field_type_18_sub_class_id <= 16'h0; // @[Control.scala 57:36]
    end else if (!(_T_1)) begin // @[Conditional.scala 40:58]
      if (!(_T_15)) begin // @[Conditional.scala 39:67]
        if (!(_T_17)) begin // @[Conditional.scala 39:67]
          classmeta_reg_desc_state_field_type_18_sub_class_id <= _GEN_755;
        end
      end
    end
    if (reset) begin // @[Control.scala 57:36]
      classmeta_reg_desc_state_field_type_18_is_host <= 1'h0; // @[Control.scala 57:36]
    end else if (!(_T_1)) begin // @[Conditional.scala 40:58]
      if (!(_T_15)) begin // @[Conditional.scala 39:67]
        if (!(_T_17)) begin // @[Conditional.scala 39:67]
          classmeta_reg_desc_state_field_type_18_is_host <= _GEN_752;
        end
      end
    end
    if (reset) begin // @[Control.scala 57:36]
      classmeta_reg_desc_state_field_type_19_is_repeated <= 1'h0; // @[Control.scala 57:36]
    end else if (!(_T_1)) begin // @[Conditional.scala 40:58]
      if (!(_T_15)) begin // @[Conditional.scala 39:67]
        if (!(_T_17)) begin // @[Conditional.scala 39:67]
          classmeta_reg_desc_state_field_type_19_is_repeated <= _GEN_757;
        end
      end
    end
    if (reset) begin // @[Control.scala 57:36]
      classmeta_reg_desc_state_field_type_19_field_type <= 5'h0; // @[Control.scala 57:36]
    end else if (!(_T_1)) begin // @[Conditional.scala 40:58]
      if (!(_T_15)) begin // @[Conditional.scala 39:67]
        if (!(_T_17)) begin // @[Conditional.scala 39:67]
          classmeta_reg_desc_state_field_type_19_field_type <= _GEN_758;
        end
      end
    end
    if (reset) begin // @[Control.scala 57:36]
      classmeta_reg_desc_state_field_type_19_sub_class_id <= 16'h0; // @[Control.scala 57:36]
    end else if (!(_T_1)) begin // @[Conditional.scala 40:58]
      if (!(_T_15)) begin // @[Conditional.scala 39:67]
        if (!(_T_17)) begin // @[Conditional.scala 39:67]
          classmeta_reg_desc_state_field_type_19_sub_class_id <= _GEN_759;
        end
      end
    end
    if (reset) begin // @[Control.scala 57:36]
      classmeta_reg_desc_state_field_type_19_is_host <= 1'h0; // @[Control.scala 57:36]
    end else if (!(_T_1)) begin // @[Conditional.scala 40:58]
      if (!(_T_15)) begin // @[Conditional.scala 39:67]
        if (!(_T_17)) begin // @[Conditional.scala 39:67]
          classmeta_reg_desc_state_field_type_19_is_host <= _GEN_756;
        end
      end
    end
    if (reset) begin // @[Control.scala 57:36]
      classmeta_reg_desc_state_field_type_20_is_repeated <= 1'h0; // @[Control.scala 57:36]
    end else if (!(_T_1)) begin // @[Conditional.scala 40:58]
      if (!(_T_15)) begin // @[Conditional.scala 39:67]
        if (!(_T_17)) begin // @[Conditional.scala 39:67]
          classmeta_reg_desc_state_field_type_20_is_repeated <= _GEN_761;
        end
      end
    end
    if (reset) begin // @[Control.scala 57:36]
      classmeta_reg_desc_state_field_type_20_field_type <= 5'h0; // @[Control.scala 57:36]
    end else if (!(_T_1)) begin // @[Conditional.scala 40:58]
      if (!(_T_15)) begin // @[Conditional.scala 39:67]
        if (!(_T_17)) begin // @[Conditional.scala 39:67]
          classmeta_reg_desc_state_field_type_20_field_type <= _GEN_762;
        end
      end
    end
    if (reset) begin // @[Control.scala 57:36]
      classmeta_reg_desc_state_field_type_20_sub_class_id <= 16'h0; // @[Control.scala 57:36]
    end else if (!(_T_1)) begin // @[Conditional.scala 40:58]
      if (!(_T_15)) begin // @[Conditional.scala 39:67]
        if (!(_T_17)) begin // @[Conditional.scala 39:67]
          classmeta_reg_desc_state_field_type_20_sub_class_id <= _GEN_763;
        end
      end
    end
    if (reset) begin // @[Control.scala 57:36]
      classmeta_reg_desc_state_field_type_20_is_host <= 1'h0; // @[Control.scala 57:36]
    end else if (!(_T_1)) begin // @[Conditional.scala 40:58]
      if (!(_T_15)) begin // @[Conditional.scala 39:67]
        if (!(_T_17)) begin // @[Conditional.scala 39:67]
          classmeta_reg_desc_state_field_type_20_is_host <= _GEN_760;
        end
      end
    end
    if (reset) begin // @[Control.scala 57:36]
      classmeta_reg_desc_state_field_type_21_is_repeated <= 1'h0; // @[Control.scala 57:36]
    end else if (!(_T_1)) begin // @[Conditional.scala 40:58]
      if (!(_T_15)) begin // @[Conditional.scala 39:67]
        if (!(_T_17)) begin // @[Conditional.scala 39:67]
          classmeta_reg_desc_state_field_type_21_is_repeated <= _GEN_765;
        end
      end
    end
    if (reset) begin // @[Control.scala 57:36]
      classmeta_reg_desc_state_field_type_21_field_type <= 5'h0; // @[Control.scala 57:36]
    end else if (!(_T_1)) begin // @[Conditional.scala 40:58]
      if (!(_T_15)) begin // @[Conditional.scala 39:67]
        if (!(_T_17)) begin // @[Conditional.scala 39:67]
          classmeta_reg_desc_state_field_type_21_field_type <= _GEN_766;
        end
      end
    end
    if (reset) begin // @[Control.scala 57:36]
      classmeta_reg_desc_state_field_type_21_sub_class_id <= 16'h0; // @[Control.scala 57:36]
    end else if (!(_T_1)) begin // @[Conditional.scala 40:58]
      if (!(_T_15)) begin // @[Conditional.scala 39:67]
        if (!(_T_17)) begin // @[Conditional.scala 39:67]
          classmeta_reg_desc_state_field_type_21_sub_class_id <= _GEN_767;
        end
      end
    end
    if (reset) begin // @[Control.scala 57:36]
      classmeta_reg_desc_state_field_type_21_is_host <= 1'h0; // @[Control.scala 57:36]
    end else if (!(_T_1)) begin // @[Conditional.scala 40:58]
      if (!(_T_15)) begin // @[Conditional.scala 39:67]
        if (!(_T_17)) begin // @[Conditional.scala 39:67]
          classmeta_reg_desc_state_field_type_21_is_host <= _GEN_764;
        end
      end
    end
    if (reset) begin // @[Control.scala 57:36]
      classmeta_reg_desc_state_field_type_22_is_repeated <= 1'h0; // @[Control.scala 57:36]
    end else if (!(_T_1)) begin // @[Conditional.scala 40:58]
      if (!(_T_15)) begin // @[Conditional.scala 39:67]
        if (!(_T_17)) begin // @[Conditional.scala 39:67]
          classmeta_reg_desc_state_field_type_22_is_repeated <= _GEN_769;
        end
      end
    end
    if (reset) begin // @[Control.scala 57:36]
      classmeta_reg_desc_state_field_type_22_field_type <= 5'h0; // @[Control.scala 57:36]
    end else if (!(_T_1)) begin // @[Conditional.scala 40:58]
      if (!(_T_15)) begin // @[Conditional.scala 39:67]
        if (!(_T_17)) begin // @[Conditional.scala 39:67]
          classmeta_reg_desc_state_field_type_22_field_type <= _GEN_770;
        end
      end
    end
    if (reset) begin // @[Control.scala 57:36]
      classmeta_reg_desc_state_field_type_22_sub_class_id <= 16'h0; // @[Control.scala 57:36]
    end else if (!(_T_1)) begin // @[Conditional.scala 40:58]
      if (!(_T_15)) begin // @[Conditional.scala 39:67]
        if (!(_T_17)) begin // @[Conditional.scala 39:67]
          classmeta_reg_desc_state_field_type_22_sub_class_id <= _GEN_771;
        end
      end
    end
    if (reset) begin // @[Control.scala 57:36]
      classmeta_reg_desc_state_field_type_22_is_host <= 1'h0; // @[Control.scala 57:36]
    end else if (!(_T_1)) begin // @[Conditional.scala 40:58]
      if (!(_T_15)) begin // @[Conditional.scala 39:67]
        if (!(_T_17)) begin // @[Conditional.scala 39:67]
          classmeta_reg_desc_state_field_type_22_is_host <= _GEN_768;
        end
      end
    end
    if (reset) begin // @[Control.scala 57:36]
      classmeta_reg_desc_state_field_type_23_is_repeated <= 1'h0; // @[Control.scala 57:36]
    end else if (!(_T_1)) begin // @[Conditional.scala 40:58]
      if (!(_T_15)) begin // @[Conditional.scala 39:67]
        if (!(_T_17)) begin // @[Conditional.scala 39:67]
          classmeta_reg_desc_state_field_type_23_is_repeated <= _GEN_773;
        end
      end
    end
    if (reset) begin // @[Control.scala 57:36]
      classmeta_reg_desc_state_field_type_23_field_type <= 5'h0; // @[Control.scala 57:36]
    end else if (!(_T_1)) begin // @[Conditional.scala 40:58]
      if (!(_T_15)) begin // @[Conditional.scala 39:67]
        if (!(_T_17)) begin // @[Conditional.scala 39:67]
          classmeta_reg_desc_state_field_type_23_field_type <= _GEN_774;
        end
      end
    end
    if (reset) begin // @[Control.scala 57:36]
      classmeta_reg_desc_state_field_type_23_sub_class_id <= 16'h0; // @[Control.scala 57:36]
    end else if (!(_T_1)) begin // @[Conditional.scala 40:58]
      if (!(_T_15)) begin // @[Conditional.scala 39:67]
        if (!(_T_17)) begin // @[Conditional.scala 39:67]
          classmeta_reg_desc_state_field_type_23_sub_class_id <= _GEN_775;
        end
      end
    end
    if (reset) begin // @[Control.scala 57:36]
      classmeta_reg_desc_state_field_type_23_is_host <= 1'h0; // @[Control.scala 57:36]
    end else if (!(_T_1)) begin // @[Conditional.scala 40:58]
      if (!(_T_15)) begin // @[Conditional.scala 39:67]
        if (!(_T_17)) begin // @[Conditional.scala 39:67]
          classmeta_reg_desc_state_field_type_23_is_host <= _GEN_772;
        end
      end
    end
    if (reset) begin // @[Control.scala 57:36]
      classmeta_reg_desc_state_field_type_24_is_repeated <= 1'h0; // @[Control.scala 57:36]
    end else if (!(_T_1)) begin // @[Conditional.scala 40:58]
      if (!(_T_15)) begin // @[Conditional.scala 39:67]
        if (!(_T_17)) begin // @[Conditional.scala 39:67]
          classmeta_reg_desc_state_field_type_24_is_repeated <= _GEN_777;
        end
      end
    end
    if (reset) begin // @[Control.scala 57:36]
      classmeta_reg_desc_state_field_type_24_field_type <= 5'h0; // @[Control.scala 57:36]
    end else if (!(_T_1)) begin // @[Conditional.scala 40:58]
      if (!(_T_15)) begin // @[Conditional.scala 39:67]
        if (!(_T_17)) begin // @[Conditional.scala 39:67]
          classmeta_reg_desc_state_field_type_24_field_type <= _GEN_778;
        end
      end
    end
    if (reset) begin // @[Control.scala 57:36]
      classmeta_reg_desc_state_field_type_24_sub_class_id <= 16'h0; // @[Control.scala 57:36]
    end else if (!(_T_1)) begin // @[Conditional.scala 40:58]
      if (!(_T_15)) begin // @[Conditional.scala 39:67]
        if (!(_T_17)) begin // @[Conditional.scala 39:67]
          classmeta_reg_desc_state_field_type_24_sub_class_id <= _GEN_779;
        end
      end
    end
    if (reset) begin // @[Control.scala 57:36]
      classmeta_reg_desc_state_field_type_24_is_host <= 1'h0; // @[Control.scala 57:36]
    end else if (!(_T_1)) begin // @[Conditional.scala 40:58]
      if (!(_T_15)) begin // @[Conditional.scala 39:67]
        if (!(_T_17)) begin // @[Conditional.scala 39:67]
          classmeta_reg_desc_state_field_type_24_is_host <= _GEN_776;
        end
      end
    end
    if (reset) begin // @[Control.scala 57:36]
      classmeta_reg_desc_state_field_type_25_is_repeated <= 1'h0; // @[Control.scala 57:36]
    end else if (!(_T_1)) begin // @[Conditional.scala 40:58]
      if (!(_T_15)) begin // @[Conditional.scala 39:67]
        if (!(_T_17)) begin // @[Conditional.scala 39:67]
          classmeta_reg_desc_state_field_type_25_is_repeated <= _GEN_781;
        end
      end
    end
    if (reset) begin // @[Control.scala 57:36]
      classmeta_reg_desc_state_field_type_25_field_type <= 5'h0; // @[Control.scala 57:36]
    end else if (!(_T_1)) begin // @[Conditional.scala 40:58]
      if (!(_T_15)) begin // @[Conditional.scala 39:67]
        if (!(_T_17)) begin // @[Conditional.scala 39:67]
          classmeta_reg_desc_state_field_type_25_field_type <= _GEN_782;
        end
      end
    end
    if (reset) begin // @[Control.scala 57:36]
      classmeta_reg_desc_state_field_type_25_sub_class_id <= 16'h0; // @[Control.scala 57:36]
    end else if (!(_T_1)) begin // @[Conditional.scala 40:58]
      if (!(_T_15)) begin // @[Conditional.scala 39:67]
        if (!(_T_17)) begin // @[Conditional.scala 39:67]
          classmeta_reg_desc_state_field_type_25_sub_class_id <= _GEN_783;
        end
      end
    end
    if (reset) begin // @[Control.scala 57:36]
      classmeta_reg_desc_state_field_type_25_is_host <= 1'h0; // @[Control.scala 57:36]
    end else if (!(_T_1)) begin // @[Conditional.scala 40:58]
      if (!(_T_15)) begin // @[Conditional.scala 39:67]
        if (!(_T_17)) begin // @[Conditional.scala 39:67]
          classmeta_reg_desc_state_field_type_25_is_host <= _GEN_780;
        end
      end
    end
    if (reset) begin // @[Control.scala 57:36]
      classmeta_reg_desc_state_field_type_26_is_repeated <= 1'h0; // @[Control.scala 57:36]
    end else if (!(_T_1)) begin // @[Conditional.scala 40:58]
      if (!(_T_15)) begin // @[Conditional.scala 39:67]
        if (!(_T_17)) begin // @[Conditional.scala 39:67]
          classmeta_reg_desc_state_field_type_26_is_repeated <= _GEN_785;
        end
      end
    end
    if (reset) begin // @[Control.scala 57:36]
      classmeta_reg_desc_state_field_type_26_field_type <= 5'h0; // @[Control.scala 57:36]
    end else if (!(_T_1)) begin // @[Conditional.scala 40:58]
      if (!(_T_15)) begin // @[Conditional.scala 39:67]
        if (!(_T_17)) begin // @[Conditional.scala 39:67]
          classmeta_reg_desc_state_field_type_26_field_type <= _GEN_786;
        end
      end
    end
    if (reset) begin // @[Control.scala 57:36]
      classmeta_reg_desc_state_field_type_26_sub_class_id <= 16'h0; // @[Control.scala 57:36]
    end else if (!(_T_1)) begin // @[Conditional.scala 40:58]
      if (!(_T_15)) begin // @[Conditional.scala 39:67]
        if (!(_T_17)) begin // @[Conditional.scala 39:67]
          classmeta_reg_desc_state_field_type_26_sub_class_id <= _GEN_787;
        end
      end
    end
    if (reset) begin // @[Control.scala 57:36]
      classmeta_reg_desc_state_field_type_26_is_host <= 1'h0; // @[Control.scala 57:36]
    end else if (!(_T_1)) begin // @[Conditional.scala 40:58]
      if (!(_T_15)) begin // @[Conditional.scala 39:67]
        if (!(_T_17)) begin // @[Conditional.scala 39:67]
          classmeta_reg_desc_state_field_type_26_is_host <= _GEN_784;
        end
      end
    end
    if (reset) begin // @[Control.scala 57:36]
      classmeta_reg_desc_state_field_type_27_is_repeated <= 1'h0; // @[Control.scala 57:36]
    end else if (!(_T_1)) begin // @[Conditional.scala 40:58]
      if (!(_T_15)) begin // @[Conditional.scala 39:67]
        if (!(_T_17)) begin // @[Conditional.scala 39:67]
          classmeta_reg_desc_state_field_type_27_is_repeated <= _GEN_789;
        end
      end
    end
    if (reset) begin // @[Control.scala 57:36]
      classmeta_reg_desc_state_field_type_27_field_type <= 5'h0; // @[Control.scala 57:36]
    end else if (!(_T_1)) begin // @[Conditional.scala 40:58]
      if (!(_T_15)) begin // @[Conditional.scala 39:67]
        if (!(_T_17)) begin // @[Conditional.scala 39:67]
          classmeta_reg_desc_state_field_type_27_field_type <= _GEN_790;
        end
      end
    end
    if (reset) begin // @[Control.scala 57:36]
      classmeta_reg_desc_state_field_type_27_sub_class_id <= 16'h0; // @[Control.scala 57:36]
    end else if (!(_T_1)) begin // @[Conditional.scala 40:58]
      if (!(_T_15)) begin // @[Conditional.scala 39:67]
        if (!(_T_17)) begin // @[Conditional.scala 39:67]
          classmeta_reg_desc_state_field_type_27_sub_class_id <= _GEN_791;
        end
      end
    end
    if (reset) begin // @[Control.scala 57:36]
      classmeta_reg_desc_state_field_type_27_is_host <= 1'h0; // @[Control.scala 57:36]
    end else if (!(_T_1)) begin // @[Conditional.scala 40:58]
      if (!(_T_15)) begin // @[Conditional.scala 39:67]
        if (!(_T_17)) begin // @[Conditional.scala 39:67]
          classmeta_reg_desc_state_field_type_27_is_host <= _GEN_788;
        end
      end
    end
    if (reset) begin // @[Control.scala 57:36]
      classmeta_reg_desc_state_field_type_28_is_repeated <= 1'h0; // @[Control.scala 57:36]
    end else if (!(_T_1)) begin // @[Conditional.scala 40:58]
      if (!(_T_15)) begin // @[Conditional.scala 39:67]
        if (!(_T_17)) begin // @[Conditional.scala 39:67]
          classmeta_reg_desc_state_field_type_28_is_repeated <= _GEN_793;
        end
      end
    end
    if (reset) begin // @[Control.scala 57:36]
      classmeta_reg_desc_state_field_type_28_field_type <= 5'h0; // @[Control.scala 57:36]
    end else if (!(_T_1)) begin // @[Conditional.scala 40:58]
      if (!(_T_15)) begin // @[Conditional.scala 39:67]
        if (!(_T_17)) begin // @[Conditional.scala 39:67]
          classmeta_reg_desc_state_field_type_28_field_type <= _GEN_794;
        end
      end
    end
    if (reset) begin // @[Control.scala 57:36]
      classmeta_reg_desc_state_field_type_28_sub_class_id <= 16'h0; // @[Control.scala 57:36]
    end else if (!(_T_1)) begin // @[Conditional.scala 40:58]
      if (!(_T_15)) begin // @[Conditional.scala 39:67]
        if (!(_T_17)) begin // @[Conditional.scala 39:67]
          classmeta_reg_desc_state_field_type_28_sub_class_id <= _GEN_795;
        end
      end
    end
    if (reset) begin // @[Control.scala 57:36]
      classmeta_reg_desc_state_field_type_28_is_host <= 1'h0; // @[Control.scala 57:36]
    end else if (!(_T_1)) begin // @[Conditional.scala 40:58]
      if (!(_T_15)) begin // @[Conditional.scala 39:67]
        if (!(_T_17)) begin // @[Conditional.scala 39:67]
          classmeta_reg_desc_state_field_type_28_is_host <= _GEN_792;
        end
      end
    end
    if (reset) begin // @[Control.scala 57:36]
      classmeta_reg_desc_state_field_type_29_is_repeated <= 1'h0; // @[Control.scala 57:36]
    end else if (!(_T_1)) begin // @[Conditional.scala 40:58]
      if (!(_T_15)) begin // @[Conditional.scala 39:67]
        if (!(_T_17)) begin // @[Conditional.scala 39:67]
          classmeta_reg_desc_state_field_type_29_is_repeated <= _GEN_797;
        end
      end
    end
    if (reset) begin // @[Control.scala 57:36]
      classmeta_reg_desc_state_field_type_29_field_type <= 5'h0; // @[Control.scala 57:36]
    end else if (!(_T_1)) begin // @[Conditional.scala 40:58]
      if (!(_T_15)) begin // @[Conditional.scala 39:67]
        if (!(_T_17)) begin // @[Conditional.scala 39:67]
          classmeta_reg_desc_state_field_type_29_field_type <= _GEN_798;
        end
      end
    end
    if (reset) begin // @[Control.scala 57:36]
      classmeta_reg_desc_state_field_type_29_sub_class_id <= 16'h0; // @[Control.scala 57:36]
    end else if (!(_T_1)) begin // @[Conditional.scala 40:58]
      if (!(_T_15)) begin // @[Conditional.scala 39:67]
        if (!(_T_17)) begin // @[Conditional.scala 39:67]
          classmeta_reg_desc_state_field_type_29_sub_class_id <= _GEN_799;
        end
      end
    end
    if (reset) begin // @[Control.scala 57:36]
      classmeta_reg_desc_state_field_type_29_is_host <= 1'h0; // @[Control.scala 57:36]
    end else if (!(_T_1)) begin // @[Conditional.scala 40:58]
      if (!(_T_15)) begin // @[Conditional.scala 39:67]
        if (!(_T_17)) begin // @[Conditional.scala 39:67]
          classmeta_reg_desc_state_field_type_29_is_host <= _GEN_796;
        end
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  s_wr = _RAND_0[2:0];
  _RAND_1 = {1{`RANDOM}};
  cur_data = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  classmeta_reg_class_id = _RAND_2[9:0];
  _RAND_3 = {1{`RANDOM}};
  classmeta_reg_desc_state_class_length = _RAND_3[15:0];
  _RAND_4 = {1{`RANDOM}};
  classmeta_reg_desc_state_max_field_num = _RAND_4[7:0];
  _RAND_5 = {1{`RANDOM}};
  classmeta_reg_desc_state_field_type_0_is_repeated = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  classmeta_reg_desc_state_field_type_0_field_type = _RAND_6[4:0];
  _RAND_7 = {1{`RANDOM}};
  classmeta_reg_desc_state_field_type_0_sub_class_id = _RAND_7[15:0];
  _RAND_8 = {1{`RANDOM}};
  classmeta_reg_desc_state_field_type_0_is_host = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  classmeta_reg_desc_state_field_type_1_is_repeated = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  classmeta_reg_desc_state_field_type_1_field_type = _RAND_10[4:0];
  _RAND_11 = {1{`RANDOM}};
  classmeta_reg_desc_state_field_type_1_sub_class_id = _RAND_11[15:0];
  _RAND_12 = {1{`RANDOM}};
  classmeta_reg_desc_state_field_type_1_is_host = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  classmeta_reg_desc_state_field_type_2_is_repeated = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  classmeta_reg_desc_state_field_type_2_field_type = _RAND_14[4:0];
  _RAND_15 = {1{`RANDOM}};
  classmeta_reg_desc_state_field_type_2_sub_class_id = _RAND_15[15:0];
  _RAND_16 = {1{`RANDOM}};
  classmeta_reg_desc_state_field_type_2_is_host = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  classmeta_reg_desc_state_field_type_3_is_repeated = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  classmeta_reg_desc_state_field_type_3_field_type = _RAND_18[4:0];
  _RAND_19 = {1{`RANDOM}};
  classmeta_reg_desc_state_field_type_3_sub_class_id = _RAND_19[15:0];
  _RAND_20 = {1{`RANDOM}};
  classmeta_reg_desc_state_field_type_3_is_host = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  classmeta_reg_desc_state_field_type_4_is_repeated = _RAND_21[0:0];
  _RAND_22 = {1{`RANDOM}};
  classmeta_reg_desc_state_field_type_4_field_type = _RAND_22[4:0];
  _RAND_23 = {1{`RANDOM}};
  classmeta_reg_desc_state_field_type_4_sub_class_id = _RAND_23[15:0];
  _RAND_24 = {1{`RANDOM}};
  classmeta_reg_desc_state_field_type_4_is_host = _RAND_24[0:0];
  _RAND_25 = {1{`RANDOM}};
  classmeta_reg_desc_state_field_type_5_is_repeated = _RAND_25[0:0];
  _RAND_26 = {1{`RANDOM}};
  classmeta_reg_desc_state_field_type_5_field_type = _RAND_26[4:0];
  _RAND_27 = {1{`RANDOM}};
  classmeta_reg_desc_state_field_type_5_sub_class_id = _RAND_27[15:0];
  _RAND_28 = {1{`RANDOM}};
  classmeta_reg_desc_state_field_type_5_is_host = _RAND_28[0:0];
  _RAND_29 = {1{`RANDOM}};
  classmeta_reg_desc_state_field_type_6_is_repeated = _RAND_29[0:0];
  _RAND_30 = {1{`RANDOM}};
  classmeta_reg_desc_state_field_type_6_field_type = _RAND_30[4:0];
  _RAND_31 = {1{`RANDOM}};
  classmeta_reg_desc_state_field_type_6_sub_class_id = _RAND_31[15:0];
  _RAND_32 = {1{`RANDOM}};
  classmeta_reg_desc_state_field_type_6_is_host = _RAND_32[0:0];
  _RAND_33 = {1{`RANDOM}};
  classmeta_reg_desc_state_field_type_7_is_repeated = _RAND_33[0:0];
  _RAND_34 = {1{`RANDOM}};
  classmeta_reg_desc_state_field_type_7_field_type = _RAND_34[4:0];
  _RAND_35 = {1{`RANDOM}};
  classmeta_reg_desc_state_field_type_7_sub_class_id = _RAND_35[15:0];
  _RAND_36 = {1{`RANDOM}};
  classmeta_reg_desc_state_field_type_7_is_host = _RAND_36[0:0];
  _RAND_37 = {1{`RANDOM}};
  classmeta_reg_desc_state_field_type_8_is_repeated = _RAND_37[0:0];
  _RAND_38 = {1{`RANDOM}};
  classmeta_reg_desc_state_field_type_8_field_type = _RAND_38[4:0];
  _RAND_39 = {1{`RANDOM}};
  classmeta_reg_desc_state_field_type_8_sub_class_id = _RAND_39[15:0];
  _RAND_40 = {1{`RANDOM}};
  classmeta_reg_desc_state_field_type_8_is_host = _RAND_40[0:0];
  _RAND_41 = {1{`RANDOM}};
  classmeta_reg_desc_state_field_type_9_is_repeated = _RAND_41[0:0];
  _RAND_42 = {1{`RANDOM}};
  classmeta_reg_desc_state_field_type_9_field_type = _RAND_42[4:0];
  _RAND_43 = {1{`RANDOM}};
  classmeta_reg_desc_state_field_type_9_sub_class_id = _RAND_43[15:0];
  _RAND_44 = {1{`RANDOM}};
  classmeta_reg_desc_state_field_type_9_is_host = _RAND_44[0:0];
  _RAND_45 = {1{`RANDOM}};
  classmeta_reg_desc_state_field_type_10_is_repeated = _RAND_45[0:0];
  _RAND_46 = {1{`RANDOM}};
  classmeta_reg_desc_state_field_type_10_field_type = _RAND_46[4:0];
  _RAND_47 = {1{`RANDOM}};
  classmeta_reg_desc_state_field_type_10_sub_class_id = _RAND_47[15:0];
  _RAND_48 = {1{`RANDOM}};
  classmeta_reg_desc_state_field_type_10_is_host = _RAND_48[0:0];
  _RAND_49 = {1{`RANDOM}};
  classmeta_reg_desc_state_field_type_11_is_repeated = _RAND_49[0:0];
  _RAND_50 = {1{`RANDOM}};
  classmeta_reg_desc_state_field_type_11_field_type = _RAND_50[4:0];
  _RAND_51 = {1{`RANDOM}};
  classmeta_reg_desc_state_field_type_11_sub_class_id = _RAND_51[15:0];
  _RAND_52 = {1{`RANDOM}};
  classmeta_reg_desc_state_field_type_11_is_host = _RAND_52[0:0];
  _RAND_53 = {1{`RANDOM}};
  classmeta_reg_desc_state_field_type_12_is_repeated = _RAND_53[0:0];
  _RAND_54 = {1{`RANDOM}};
  classmeta_reg_desc_state_field_type_12_field_type = _RAND_54[4:0];
  _RAND_55 = {1{`RANDOM}};
  classmeta_reg_desc_state_field_type_12_sub_class_id = _RAND_55[15:0];
  _RAND_56 = {1{`RANDOM}};
  classmeta_reg_desc_state_field_type_12_is_host = _RAND_56[0:0];
  _RAND_57 = {1{`RANDOM}};
  classmeta_reg_desc_state_field_type_13_is_repeated = _RAND_57[0:0];
  _RAND_58 = {1{`RANDOM}};
  classmeta_reg_desc_state_field_type_13_field_type = _RAND_58[4:0];
  _RAND_59 = {1{`RANDOM}};
  classmeta_reg_desc_state_field_type_13_sub_class_id = _RAND_59[15:0];
  _RAND_60 = {1{`RANDOM}};
  classmeta_reg_desc_state_field_type_13_is_host = _RAND_60[0:0];
  _RAND_61 = {1{`RANDOM}};
  classmeta_reg_desc_state_field_type_14_is_repeated = _RAND_61[0:0];
  _RAND_62 = {1{`RANDOM}};
  classmeta_reg_desc_state_field_type_14_field_type = _RAND_62[4:0];
  _RAND_63 = {1{`RANDOM}};
  classmeta_reg_desc_state_field_type_14_sub_class_id = _RAND_63[15:0];
  _RAND_64 = {1{`RANDOM}};
  classmeta_reg_desc_state_field_type_14_is_host = _RAND_64[0:0];
  _RAND_65 = {1{`RANDOM}};
  classmeta_reg_desc_state_field_type_15_is_repeated = _RAND_65[0:0];
  _RAND_66 = {1{`RANDOM}};
  classmeta_reg_desc_state_field_type_15_field_type = _RAND_66[4:0];
  _RAND_67 = {1{`RANDOM}};
  classmeta_reg_desc_state_field_type_15_sub_class_id = _RAND_67[15:0];
  _RAND_68 = {1{`RANDOM}};
  classmeta_reg_desc_state_field_type_15_is_host = _RAND_68[0:0];
  _RAND_69 = {1{`RANDOM}};
  classmeta_reg_desc_state_field_type_16_is_repeated = _RAND_69[0:0];
  _RAND_70 = {1{`RANDOM}};
  classmeta_reg_desc_state_field_type_16_field_type = _RAND_70[4:0];
  _RAND_71 = {1{`RANDOM}};
  classmeta_reg_desc_state_field_type_16_sub_class_id = _RAND_71[15:0];
  _RAND_72 = {1{`RANDOM}};
  classmeta_reg_desc_state_field_type_16_is_host = _RAND_72[0:0];
  _RAND_73 = {1{`RANDOM}};
  classmeta_reg_desc_state_field_type_17_is_repeated = _RAND_73[0:0];
  _RAND_74 = {1{`RANDOM}};
  classmeta_reg_desc_state_field_type_17_field_type = _RAND_74[4:0];
  _RAND_75 = {1{`RANDOM}};
  classmeta_reg_desc_state_field_type_17_sub_class_id = _RAND_75[15:0];
  _RAND_76 = {1{`RANDOM}};
  classmeta_reg_desc_state_field_type_17_is_host = _RAND_76[0:0];
  _RAND_77 = {1{`RANDOM}};
  classmeta_reg_desc_state_field_type_18_is_repeated = _RAND_77[0:0];
  _RAND_78 = {1{`RANDOM}};
  classmeta_reg_desc_state_field_type_18_field_type = _RAND_78[4:0];
  _RAND_79 = {1{`RANDOM}};
  classmeta_reg_desc_state_field_type_18_sub_class_id = _RAND_79[15:0];
  _RAND_80 = {1{`RANDOM}};
  classmeta_reg_desc_state_field_type_18_is_host = _RAND_80[0:0];
  _RAND_81 = {1{`RANDOM}};
  classmeta_reg_desc_state_field_type_19_is_repeated = _RAND_81[0:0];
  _RAND_82 = {1{`RANDOM}};
  classmeta_reg_desc_state_field_type_19_field_type = _RAND_82[4:0];
  _RAND_83 = {1{`RANDOM}};
  classmeta_reg_desc_state_field_type_19_sub_class_id = _RAND_83[15:0];
  _RAND_84 = {1{`RANDOM}};
  classmeta_reg_desc_state_field_type_19_is_host = _RAND_84[0:0];
  _RAND_85 = {1{`RANDOM}};
  classmeta_reg_desc_state_field_type_20_is_repeated = _RAND_85[0:0];
  _RAND_86 = {1{`RANDOM}};
  classmeta_reg_desc_state_field_type_20_field_type = _RAND_86[4:0];
  _RAND_87 = {1{`RANDOM}};
  classmeta_reg_desc_state_field_type_20_sub_class_id = _RAND_87[15:0];
  _RAND_88 = {1{`RANDOM}};
  classmeta_reg_desc_state_field_type_20_is_host = _RAND_88[0:0];
  _RAND_89 = {1{`RANDOM}};
  classmeta_reg_desc_state_field_type_21_is_repeated = _RAND_89[0:0];
  _RAND_90 = {1{`RANDOM}};
  classmeta_reg_desc_state_field_type_21_field_type = _RAND_90[4:0];
  _RAND_91 = {1{`RANDOM}};
  classmeta_reg_desc_state_field_type_21_sub_class_id = _RAND_91[15:0];
  _RAND_92 = {1{`RANDOM}};
  classmeta_reg_desc_state_field_type_21_is_host = _RAND_92[0:0];
  _RAND_93 = {1{`RANDOM}};
  classmeta_reg_desc_state_field_type_22_is_repeated = _RAND_93[0:0];
  _RAND_94 = {1{`RANDOM}};
  classmeta_reg_desc_state_field_type_22_field_type = _RAND_94[4:0];
  _RAND_95 = {1{`RANDOM}};
  classmeta_reg_desc_state_field_type_22_sub_class_id = _RAND_95[15:0];
  _RAND_96 = {1{`RANDOM}};
  classmeta_reg_desc_state_field_type_22_is_host = _RAND_96[0:0];
  _RAND_97 = {1{`RANDOM}};
  classmeta_reg_desc_state_field_type_23_is_repeated = _RAND_97[0:0];
  _RAND_98 = {1{`RANDOM}};
  classmeta_reg_desc_state_field_type_23_field_type = _RAND_98[4:0];
  _RAND_99 = {1{`RANDOM}};
  classmeta_reg_desc_state_field_type_23_sub_class_id = _RAND_99[15:0];
  _RAND_100 = {1{`RANDOM}};
  classmeta_reg_desc_state_field_type_23_is_host = _RAND_100[0:0];
  _RAND_101 = {1{`RANDOM}};
  classmeta_reg_desc_state_field_type_24_is_repeated = _RAND_101[0:0];
  _RAND_102 = {1{`RANDOM}};
  classmeta_reg_desc_state_field_type_24_field_type = _RAND_102[4:0];
  _RAND_103 = {1{`RANDOM}};
  classmeta_reg_desc_state_field_type_24_sub_class_id = _RAND_103[15:0];
  _RAND_104 = {1{`RANDOM}};
  classmeta_reg_desc_state_field_type_24_is_host = _RAND_104[0:0];
  _RAND_105 = {1{`RANDOM}};
  classmeta_reg_desc_state_field_type_25_is_repeated = _RAND_105[0:0];
  _RAND_106 = {1{`RANDOM}};
  classmeta_reg_desc_state_field_type_25_field_type = _RAND_106[4:0];
  _RAND_107 = {1{`RANDOM}};
  classmeta_reg_desc_state_field_type_25_sub_class_id = _RAND_107[15:0];
  _RAND_108 = {1{`RANDOM}};
  classmeta_reg_desc_state_field_type_25_is_host = _RAND_108[0:0];
  _RAND_109 = {1{`RANDOM}};
  classmeta_reg_desc_state_field_type_26_is_repeated = _RAND_109[0:0];
  _RAND_110 = {1{`RANDOM}};
  classmeta_reg_desc_state_field_type_26_field_type = _RAND_110[4:0];
  _RAND_111 = {1{`RANDOM}};
  classmeta_reg_desc_state_field_type_26_sub_class_id = _RAND_111[15:0];
  _RAND_112 = {1{`RANDOM}};
  classmeta_reg_desc_state_field_type_26_is_host = _RAND_112[0:0];
  _RAND_113 = {1{`RANDOM}};
  classmeta_reg_desc_state_field_type_27_is_repeated = _RAND_113[0:0];
  _RAND_114 = {1{`RANDOM}};
  classmeta_reg_desc_state_field_type_27_field_type = _RAND_114[4:0];
  _RAND_115 = {1{`RANDOM}};
  classmeta_reg_desc_state_field_type_27_sub_class_id = _RAND_115[15:0];
  _RAND_116 = {1{`RANDOM}};
  classmeta_reg_desc_state_field_type_27_is_host = _RAND_116[0:0];
  _RAND_117 = {1{`RANDOM}};
  classmeta_reg_desc_state_field_type_28_is_repeated = _RAND_117[0:0];
  _RAND_118 = {1{`RANDOM}};
  classmeta_reg_desc_state_field_type_28_field_type = _RAND_118[4:0];
  _RAND_119 = {1{`RANDOM}};
  classmeta_reg_desc_state_field_type_28_sub_class_id = _RAND_119[15:0];
  _RAND_120 = {1{`RANDOM}};
  classmeta_reg_desc_state_field_type_28_is_host = _RAND_120[0:0];
  _RAND_121 = {1{`RANDOM}};
  classmeta_reg_desc_state_field_type_29_is_repeated = _RAND_121[0:0];
  _RAND_122 = {1{`RANDOM}};
  classmeta_reg_desc_state_field_type_29_field_type = _RAND_122[4:0];
  _RAND_123 = {1{`RANDOM}};
  classmeta_reg_desc_state_field_type_29_sub_class_id = _RAND_123[15:0];
  _RAND_124 = {1{`RANDOM}};
  classmeta_reg_desc_state_field_type_29_is_host = _RAND_124[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module AlveoDynamicTop(
  input          clock,
  input          reset,
  input          io_sysClk,
  input          io_serClk,
  input          io_cmacClk,
  output [3:0]   io_cmacPin_tx_p,
  output [3:0]   io_cmacPin_tx_n,
  input  [3:0]   io_cmacPin_rx_p,
  input  [3:0]   io_cmacPin_rx_n,
  input          io_cmacPin_gt_clk_p,
  input          io_cmacPin_gt_clk_n,
  output [3:0]   io_cmacPin2_tx_p,
  output [3:0]   io_cmacPin2_tx_n,
  input  [3:0]   io_cmacPin2_rx_p,
  input  [3:0]   io_cmacPin2_rx_n,
  input          io_cmacPin2_gt_clk_p,
  input          io_cmacPin2_gt_clk_n,
  input          io_ddrPort2_clk,
  input          io_ddrPort2_rst,
  input          io_ddrPort2_axi_aw_ready,
  output         io_ddrPort2_axi_aw_valid,
  output [33:0]  io_ddrPort2_axi_aw_bits_addr,
  output [1:0]   io_ddrPort2_axi_aw_bits_burst,
  output [3:0]   io_ddrPort2_axi_aw_bits_cache,
  output [3:0]   io_ddrPort2_axi_aw_bits_id,
  output [7:0]   io_ddrPort2_axi_aw_bits_len,
  output         io_ddrPort2_axi_aw_bits_lock,
  output [2:0]   io_ddrPort2_axi_aw_bits_prot,
  output [3:0]   io_ddrPort2_axi_aw_bits_qos,
  output [3:0]   io_ddrPort2_axi_aw_bits_region,
  output [2:0]   io_ddrPort2_axi_aw_bits_size,
  input          io_ddrPort2_axi_ar_ready,
  output         io_ddrPort2_axi_ar_valid,
  output [33:0]  io_ddrPort2_axi_ar_bits_addr,
  output [1:0]   io_ddrPort2_axi_ar_bits_burst,
  output [3:0]   io_ddrPort2_axi_ar_bits_cache,
  output [3:0]   io_ddrPort2_axi_ar_bits_id,
  output [7:0]   io_ddrPort2_axi_ar_bits_len,
  output         io_ddrPort2_axi_ar_bits_lock,
  output [2:0]   io_ddrPort2_axi_ar_bits_prot,
  output [3:0]   io_ddrPort2_axi_ar_bits_qos,
  output [3:0]   io_ddrPort2_axi_ar_bits_region,
  output [2:0]   io_ddrPort2_axi_ar_bits_size,
  input          io_ddrPort2_axi_w_ready,
  output         io_ddrPort2_axi_w_valid,
  output [511:0] io_ddrPort2_axi_w_bits_data,
  output         io_ddrPort2_axi_w_bits_last,
  output [63:0]  io_ddrPort2_axi_w_bits_strb,
  output         io_ddrPort2_axi_r_ready,
  input          io_ddrPort2_axi_r_valid,
  input  [511:0] io_ddrPort2_axi_r_bits_data,
  input          io_ddrPort2_axi_r_bits_last,
  input  [1:0]   io_ddrPort2_axi_r_bits_resp,
  input  [3:0]   io_ddrPort2_axi_r_bits_id,
  output         io_ddrPort2_axi_b_ready,
  input          io_ddrPort2_axi_b_valid,
  input  [3:0]   io_ddrPort2_axi_b_bits_id,
  input  [1:0]   io_ddrPort2_axi_b_bits_resp,
  input          io_qdma_axi_aclk,
  input          io_qdma_axi_aresetn,
  input  [3:0]   io_qdma_m_axib_awid,
  input  [63:0]  io_qdma_m_axib_awaddr,
  input  [7:0]   io_qdma_m_axib_awlen,
  input  [2:0]   io_qdma_m_axib_awsize,
  input  [1:0]   io_qdma_m_axib_awburst,
  input  [2:0]   io_qdma_m_axib_awprot,
  input          io_qdma_m_axib_awlock,
  input  [3:0]   io_qdma_m_axib_awcache,
  input          io_qdma_m_axib_awvalid,
  output         io_qdma_m_axib_awready,
  input  [511:0] io_qdma_m_axib_wdata,
  input  [63:0]  io_qdma_m_axib_wstrb,
  input          io_qdma_m_axib_wlast,
  input          io_qdma_m_axib_wvalid,
  output         io_qdma_m_axib_wready,
  output [3:0]   io_qdma_m_axib_bid,
  output [1:0]   io_qdma_m_axib_bresp,
  output         io_qdma_m_axib_bvalid,
  input          io_qdma_m_axib_bready,
  input  [3:0]   io_qdma_m_axib_arid,
  input  [63:0]  io_qdma_m_axib_araddr,
  input  [7:0]   io_qdma_m_axib_arlen,
  input  [2:0]   io_qdma_m_axib_arsize,
  input  [1:0]   io_qdma_m_axib_arburst,
  input  [2:0]   io_qdma_m_axib_arprot,
  input          io_qdma_m_axib_arlock,
  input  [3:0]   io_qdma_m_axib_arcache,
  input          io_qdma_m_axib_arvalid,
  output         io_qdma_m_axib_arready,
  output [3:0]   io_qdma_m_axib_rid,
  output [511:0] io_qdma_m_axib_rdata,
  output [1:0]   io_qdma_m_axib_rresp,
  output         io_qdma_m_axib_rlast,
  output         io_qdma_m_axib_rvalid,
  input          io_qdma_m_axib_rready,
  input  [31:0]  io_qdma_m_axil_awaddr,
  input          io_qdma_m_axil_awvalid,
  output         io_qdma_m_axil_awready,
  input  [31:0]  io_qdma_m_axil_wdata,
  input  [3:0]   io_qdma_m_axil_wstrb,
  input          io_qdma_m_axil_wvalid,
  output         io_qdma_m_axil_wready,
  output [1:0]   io_qdma_m_axil_bresp,
  output         io_qdma_m_axil_bvalid,
  input          io_qdma_m_axil_bready,
  input  [31:0]  io_qdma_m_axil_araddr,
  input          io_qdma_m_axil_arvalid,
  output         io_qdma_m_axil_arready,
  output [31:0]  io_qdma_m_axil_rdata,
  output [1:0]   io_qdma_m_axil_rresp,
  output         io_qdma_m_axil_rvalid,
  input          io_qdma_m_axil_rready,
  output         io_qdma_soft_reset_n,
  output [63:0]  io_qdma_h2c_byp_in_st_addr,
  output [31:0]  io_qdma_h2c_byp_in_st_len,
  output         io_qdma_h2c_byp_in_st_eop,
  output         io_qdma_h2c_byp_in_st_sop,
  output         io_qdma_h2c_byp_in_st_mrkr_req,
  output         io_qdma_h2c_byp_in_st_sdi,
  output [10:0]  io_qdma_h2c_byp_in_st_qid,
  output         io_qdma_h2c_byp_in_st_error,
  output [7:0]   io_qdma_h2c_byp_in_st_func,
  output [15:0]  io_qdma_h2c_byp_in_st_cidx,
  output [2:0]   io_qdma_h2c_byp_in_st_port_id,
  output         io_qdma_h2c_byp_in_st_no_dma,
  output         io_qdma_h2c_byp_in_st_vld,
  input          io_qdma_h2c_byp_in_st_rdy,
  output [63:0]  io_qdma_c2h_byp_in_st_csh_addr,
  output [10:0]  io_qdma_c2h_byp_in_st_csh_qid,
  output         io_qdma_c2h_byp_in_st_csh_error,
  output [7:0]   io_qdma_c2h_byp_in_st_csh_func,
  output [2:0]   io_qdma_c2h_byp_in_st_csh_port_id,
  output [6:0]   io_qdma_c2h_byp_in_st_csh_pfch_tag,
  output         io_qdma_c2h_byp_in_st_csh_vld,
  input          io_qdma_c2h_byp_in_st_csh_rdy,
  output [511:0] io_qdma_s_axis_c2h_tdata,
  output [31:0]  io_qdma_s_axis_c2h_tcrc,
  output         io_qdma_s_axis_c2h_ctrl_marker,
  output [6:0]   io_qdma_s_axis_c2h_ctrl_ecc,
  output [31:0]  io_qdma_s_axis_c2h_ctrl_len,
  output [2:0]   io_qdma_s_axis_c2h_ctrl_port_id,
  output [10:0]  io_qdma_s_axis_c2h_ctrl_qid,
  output         io_qdma_s_axis_c2h_ctrl_has_cmpt,
  output [5:0]   io_qdma_s_axis_c2h_mty,
  output         io_qdma_s_axis_c2h_tlast,
  output         io_qdma_s_axis_c2h_tvalid,
  input          io_qdma_s_axis_c2h_tready,
  input  [511:0] io_qdma_m_axis_h2c_tdata,
  input  [31:0]  io_qdma_m_axis_h2c_tcrc,
  input  [10:0]  io_qdma_m_axis_h2c_tuser_qid,
  input  [2:0]   io_qdma_m_axis_h2c_tuser_port_id,
  input          io_qdma_m_axis_h2c_tuser_err,
  input  [31:0]  io_qdma_m_axis_h2c_tuser_mdata,
  input  [5:0]   io_qdma_m_axis_h2c_tuser_mty,
  input          io_qdma_m_axis_h2c_tuser_zero_byte,
  input          io_qdma_m_axis_h2c_tlast,
  input          io_qdma_m_axis_h2c_tvalid,
  output         io_qdma_m_axis_h2c_tready,
  input          io_qdma_axis_c2h_status_drop,
  input          io_qdma_axis_c2h_status_last,
  input          io_qdma_axis_c2h_status_cmp,
  input          io_qdma_axis_c2h_status_valid,
  input  [10:0]  io_qdma_axis_c2h_status_qid,
  output [511:0] io_qdma_s_axis_c2h_cmpt_tdata,
  output [1:0]   io_qdma_s_axis_c2h_cmpt_size,
  output [15:0]  io_qdma_s_axis_c2h_cmpt_dpar,
  output         io_qdma_s_axis_c2h_cmpt_tvalid,
  input          io_qdma_s_axis_c2h_cmpt_tready,
  output [10:0]  io_qdma_s_axis_c2h_cmpt_ctrl_qid,
  output [1:0]   io_qdma_s_axis_c2h_cmpt_ctrl_cmpt_type,
  output [15:0]  io_qdma_s_axis_c2h_cmpt_ctrl_wait_pld_pkt_id,
  output         io_qdma_s_axis_c2h_cmpt_ctrl_no_wrb_marker,
  output [2:0]   io_qdma_s_axis_c2h_cmpt_ctrl_port_id,
  output         io_qdma_s_axis_c2h_cmpt_ctrl_marker,
  output         io_qdma_s_axis_c2h_cmpt_ctrl_user_trig,
  output [2:0]   io_qdma_s_axis_c2h_cmpt_ctrl_col_idx,
  output [2:0]   io_qdma_s_axis_c2h_cmpt_ctrl_err_idx,
  output         io_qdma_h2c_byp_out_rdy,
  output         io_qdma_c2h_byp_out_rdy,
  output         io_qdma_tm_dsc_sts_rdy,
  output         io_qdma_dsc_crdt_in_vld,
  input          io_qdma_dsc_crdt_in_rdy,
  output         io_qdma_dsc_crdt_in_dir,
  output         io_qdma_dsc_crdt_in_fence,
  output [10:0]  io_qdma_dsc_crdt_in_qid,
  output [15:0]  io_qdma_dsc_crdt_in_crdt,
  output         io_qdma_qsts_out_rdy,
  output         io_qdma_usr_irq_in_vld,
  output [10:0]  io_qdma_usr_irq_in_vec,
  output [7:0]   io_qdma_usr_irq_in_fnc,
  input          io_qdma_usr_irq_out_ack,
  input          io_qdma_usr_irq_out_fail,
  input          S_BSCAN_drck,
  input          S_BSCAN_shift,
  input          S_BSCAN_tdi,
  input          S_BSCAN_update,
  input          S_BSCAN_sel,
  output         S_BSCAN_tdo,
  input          S_BSCAN_tms,
  input          S_BSCAN_tck,
  input          S_BSCAN_runtest,
  input          S_BSCAN_reset,
  input          S_BSCAN_capture,
  input          S_BSCAN_bscanid_en
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
`endif // RANDOMIZE_REG_INIT
  wire  dbgBridgeInst_clk; // @[DebugBridge.scala 58:37]
  wire  dbgBridgeInst_S_BSCAN_drck; // @[DebugBridge.scala 58:37]
  wire  dbgBridgeInst_S_BSCAN_shift; // @[DebugBridge.scala 58:37]
  wire  dbgBridgeInst_S_BSCAN_tdi; // @[DebugBridge.scala 58:37]
  wire  dbgBridgeInst_S_BSCAN_update; // @[DebugBridge.scala 58:37]
  wire  dbgBridgeInst_S_BSCAN_sel; // @[DebugBridge.scala 58:37]
  wire  dbgBridgeInst_S_BSCAN_tdo; // @[DebugBridge.scala 58:37]
  wire  dbgBridgeInst_S_BSCAN_tms; // @[DebugBridge.scala 58:37]
  wire  dbgBridgeInst_S_BSCAN_tck; // @[DebugBridge.scala 58:37]
  wire  dbgBridgeInst_S_BSCAN_runtest; // @[DebugBridge.scala 58:37]
  wire  dbgBridgeInst_S_BSCAN_reset; // @[DebugBridge.scala 58:37]
  wire  dbgBridgeInst_S_BSCAN_capture; // @[DebugBridge.scala 58:37]
  wire  dbgBridgeInst_S_BSCAN_bscanid_en; // @[DebugBridge.scala 58:37]
  wire  hbmDriver_clock; // @[FpgaCloudSerHw.scala 49:70]
  wire  hbmDriver_io_hbm_clk; // @[FpgaCloudSerHw.scala 49:70]
  wire  hbmDriver_io_hbm_rstn; // @[FpgaCloudSerHw.scala 49:70]
  wire  qdma_io_qdma_port_axi_aclk; // @[FpgaCloudSerHw.scala 68:26]
  wire  qdma_io_qdma_port_axi_aresetn; // @[FpgaCloudSerHw.scala 68:26]
  wire [3:0] qdma_io_qdma_port_m_axib_awid; // @[FpgaCloudSerHw.scala 68:26]
  wire [63:0] qdma_io_qdma_port_m_axib_awaddr; // @[FpgaCloudSerHw.scala 68:26]
  wire [7:0] qdma_io_qdma_port_m_axib_awlen; // @[FpgaCloudSerHw.scala 68:26]
  wire [2:0] qdma_io_qdma_port_m_axib_awsize; // @[FpgaCloudSerHw.scala 68:26]
  wire [1:0] qdma_io_qdma_port_m_axib_awburst; // @[FpgaCloudSerHw.scala 68:26]
  wire [2:0] qdma_io_qdma_port_m_axib_awprot; // @[FpgaCloudSerHw.scala 68:26]
  wire  qdma_io_qdma_port_m_axib_awlock; // @[FpgaCloudSerHw.scala 68:26]
  wire [3:0] qdma_io_qdma_port_m_axib_awcache; // @[FpgaCloudSerHw.scala 68:26]
  wire  qdma_io_qdma_port_m_axib_awvalid; // @[FpgaCloudSerHw.scala 68:26]
  wire  qdma_io_qdma_port_m_axib_awready; // @[FpgaCloudSerHw.scala 68:26]
  wire [511:0] qdma_io_qdma_port_m_axib_wdata; // @[FpgaCloudSerHw.scala 68:26]
  wire [63:0] qdma_io_qdma_port_m_axib_wstrb; // @[FpgaCloudSerHw.scala 68:26]
  wire  qdma_io_qdma_port_m_axib_wlast; // @[FpgaCloudSerHw.scala 68:26]
  wire  qdma_io_qdma_port_m_axib_wvalid; // @[FpgaCloudSerHw.scala 68:26]
  wire  qdma_io_qdma_port_m_axib_wready; // @[FpgaCloudSerHw.scala 68:26]
  wire [3:0] qdma_io_qdma_port_m_axib_bid; // @[FpgaCloudSerHw.scala 68:26]
  wire [1:0] qdma_io_qdma_port_m_axib_bresp; // @[FpgaCloudSerHw.scala 68:26]
  wire  qdma_io_qdma_port_m_axib_bvalid; // @[FpgaCloudSerHw.scala 68:26]
  wire  qdma_io_qdma_port_m_axib_bready; // @[FpgaCloudSerHw.scala 68:26]
  wire [3:0] qdma_io_qdma_port_m_axib_arid; // @[FpgaCloudSerHw.scala 68:26]
  wire [63:0] qdma_io_qdma_port_m_axib_araddr; // @[FpgaCloudSerHw.scala 68:26]
  wire [7:0] qdma_io_qdma_port_m_axib_arlen; // @[FpgaCloudSerHw.scala 68:26]
  wire [2:0] qdma_io_qdma_port_m_axib_arsize; // @[FpgaCloudSerHw.scala 68:26]
  wire [1:0] qdma_io_qdma_port_m_axib_arburst; // @[FpgaCloudSerHw.scala 68:26]
  wire [2:0] qdma_io_qdma_port_m_axib_arprot; // @[FpgaCloudSerHw.scala 68:26]
  wire  qdma_io_qdma_port_m_axib_arlock; // @[FpgaCloudSerHw.scala 68:26]
  wire [3:0] qdma_io_qdma_port_m_axib_arcache; // @[FpgaCloudSerHw.scala 68:26]
  wire  qdma_io_qdma_port_m_axib_arvalid; // @[FpgaCloudSerHw.scala 68:26]
  wire  qdma_io_qdma_port_m_axib_arready; // @[FpgaCloudSerHw.scala 68:26]
  wire [3:0] qdma_io_qdma_port_m_axib_rid; // @[FpgaCloudSerHw.scala 68:26]
  wire [511:0] qdma_io_qdma_port_m_axib_rdata; // @[FpgaCloudSerHw.scala 68:26]
  wire [1:0] qdma_io_qdma_port_m_axib_rresp; // @[FpgaCloudSerHw.scala 68:26]
  wire  qdma_io_qdma_port_m_axib_rlast; // @[FpgaCloudSerHw.scala 68:26]
  wire  qdma_io_qdma_port_m_axib_rvalid; // @[FpgaCloudSerHw.scala 68:26]
  wire  qdma_io_qdma_port_m_axib_rready; // @[FpgaCloudSerHw.scala 68:26]
  wire [31:0] qdma_io_qdma_port_m_axil_awaddr; // @[FpgaCloudSerHw.scala 68:26]
  wire  qdma_io_qdma_port_m_axil_awvalid; // @[FpgaCloudSerHw.scala 68:26]
  wire  qdma_io_qdma_port_m_axil_awready; // @[FpgaCloudSerHw.scala 68:26]
  wire [31:0] qdma_io_qdma_port_m_axil_wdata; // @[FpgaCloudSerHw.scala 68:26]
  wire [3:0] qdma_io_qdma_port_m_axil_wstrb; // @[FpgaCloudSerHw.scala 68:26]
  wire  qdma_io_qdma_port_m_axil_wvalid; // @[FpgaCloudSerHw.scala 68:26]
  wire  qdma_io_qdma_port_m_axil_wready; // @[FpgaCloudSerHw.scala 68:26]
  wire [1:0] qdma_io_qdma_port_m_axil_bresp; // @[FpgaCloudSerHw.scala 68:26]
  wire  qdma_io_qdma_port_m_axil_bvalid; // @[FpgaCloudSerHw.scala 68:26]
  wire  qdma_io_qdma_port_m_axil_bready; // @[FpgaCloudSerHw.scala 68:26]
  wire [31:0] qdma_io_qdma_port_m_axil_araddr; // @[FpgaCloudSerHw.scala 68:26]
  wire  qdma_io_qdma_port_m_axil_arvalid; // @[FpgaCloudSerHw.scala 68:26]
  wire  qdma_io_qdma_port_m_axil_arready; // @[FpgaCloudSerHw.scala 68:26]
  wire [31:0] qdma_io_qdma_port_m_axil_rdata; // @[FpgaCloudSerHw.scala 68:26]
  wire [1:0] qdma_io_qdma_port_m_axil_rresp; // @[FpgaCloudSerHw.scala 68:26]
  wire  qdma_io_qdma_port_m_axil_rvalid; // @[FpgaCloudSerHw.scala 68:26]
  wire  qdma_io_qdma_port_m_axil_rready; // @[FpgaCloudSerHw.scala 68:26]
  wire [63:0] qdma_io_qdma_port_h2c_byp_in_st_addr; // @[FpgaCloudSerHw.scala 68:26]
  wire [31:0] qdma_io_qdma_port_h2c_byp_in_st_len; // @[FpgaCloudSerHw.scala 68:26]
  wire  qdma_io_qdma_port_h2c_byp_in_st_eop; // @[FpgaCloudSerHw.scala 68:26]
  wire  qdma_io_qdma_port_h2c_byp_in_st_sop; // @[FpgaCloudSerHw.scala 68:26]
  wire  qdma_io_qdma_port_h2c_byp_in_st_mrkr_req; // @[FpgaCloudSerHw.scala 68:26]
  wire  qdma_io_qdma_port_h2c_byp_in_st_sdi; // @[FpgaCloudSerHw.scala 68:26]
  wire [10:0] qdma_io_qdma_port_h2c_byp_in_st_qid; // @[FpgaCloudSerHw.scala 68:26]
  wire  qdma_io_qdma_port_h2c_byp_in_st_error; // @[FpgaCloudSerHw.scala 68:26]
  wire [7:0] qdma_io_qdma_port_h2c_byp_in_st_func; // @[FpgaCloudSerHw.scala 68:26]
  wire [15:0] qdma_io_qdma_port_h2c_byp_in_st_cidx; // @[FpgaCloudSerHw.scala 68:26]
  wire [2:0] qdma_io_qdma_port_h2c_byp_in_st_port_id; // @[FpgaCloudSerHw.scala 68:26]
  wire  qdma_io_qdma_port_h2c_byp_in_st_no_dma; // @[FpgaCloudSerHw.scala 68:26]
  wire  qdma_io_qdma_port_h2c_byp_in_st_vld; // @[FpgaCloudSerHw.scala 68:26]
  wire  qdma_io_qdma_port_h2c_byp_in_st_rdy; // @[FpgaCloudSerHw.scala 68:26]
  wire [63:0] qdma_io_qdma_port_c2h_byp_in_st_csh_addr; // @[FpgaCloudSerHw.scala 68:26]
  wire [10:0] qdma_io_qdma_port_c2h_byp_in_st_csh_qid; // @[FpgaCloudSerHw.scala 68:26]
  wire  qdma_io_qdma_port_c2h_byp_in_st_csh_error; // @[FpgaCloudSerHw.scala 68:26]
  wire [7:0] qdma_io_qdma_port_c2h_byp_in_st_csh_func; // @[FpgaCloudSerHw.scala 68:26]
  wire [2:0] qdma_io_qdma_port_c2h_byp_in_st_csh_port_id; // @[FpgaCloudSerHw.scala 68:26]
  wire [6:0] qdma_io_qdma_port_c2h_byp_in_st_csh_pfch_tag; // @[FpgaCloudSerHw.scala 68:26]
  wire  qdma_io_qdma_port_c2h_byp_in_st_csh_vld; // @[FpgaCloudSerHw.scala 68:26]
  wire  qdma_io_qdma_port_c2h_byp_in_st_csh_rdy; // @[FpgaCloudSerHw.scala 68:26]
  wire [511:0] qdma_io_qdma_port_s_axis_c2h_tdata; // @[FpgaCloudSerHw.scala 68:26]
  wire [31:0] qdma_io_qdma_port_s_axis_c2h_tcrc; // @[FpgaCloudSerHw.scala 68:26]
  wire  qdma_io_qdma_port_s_axis_c2h_ctrl_marker; // @[FpgaCloudSerHw.scala 68:26]
  wire [6:0] qdma_io_qdma_port_s_axis_c2h_ctrl_ecc; // @[FpgaCloudSerHw.scala 68:26]
  wire [31:0] qdma_io_qdma_port_s_axis_c2h_ctrl_len; // @[FpgaCloudSerHw.scala 68:26]
  wire [2:0] qdma_io_qdma_port_s_axis_c2h_ctrl_port_id; // @[FpgaCloudSerHw.scala 68:26]
  wire [10:0] qdma_io_qdma_port_s_axis_c2h_ctrl_qid; // @[FpgaCloudSerHw.scala 68:26]
  wire  qdma_io_qdma_port_s_axis_c2h_ctrl_has_cmpt; // @[FpgaCloudSerHw.scala 68:26]
  wire [5:0] qdma_io_qdma_port_s_axis_c2h_mty; // @[FpgaCloudSerHw.scala 68:26]
  wire  qdma_io_qdma_port_s_axis_c2h_tlast; // @[FpgaCloudSerHw.scala 68:26]
  wire  qdma_io_qdma_port_s_axis_c2h_tvalid; // @[FpgaCloudSerHw.scala 68:26]
  wire  qdma_io_qdma_port_s_axis_c2h_tready; // @[FpgaCloudSerHw.scala 68:26]
  wire [511:0] qdma_io_qdma_port_m_axis_h2c_tdata; // @[FpgaCloudSerHw.scala 68:26]
  wire [31:0] qdma_io_qdma_port_m_axis_h2c_tcrc; // @[FpgaCloudSerHw.scala 68:26]
  wire [10:0] qdma_io_qdma_port_m_axis_h2c_tuser_qid; // @[FpgaCloudSerHw.scala 68:26]
  wire [2:0] qdma_io_qdma_port_m_axis_h2c_tuser_port_id; // @[FpgaCloudSerHw.scala 68:26]
  wire  qdma_io_qdma_port_m_axis_h2c_tuser_err; // @[FpgaCloudSerHw.scala 68:26]
  wire [31:0] qdma_io_qdma_port_m_axis_h2c_tuser_mdata; // @[FpgaCloudSerHw.scala 68:26]
  wire [5:0] qdma_io_qdma_port_m_axis_h2c_tuser_mty; // @[FpgaCloudSerHw.scala 68:26]
  wire  qdma_io_qdma_port_m_axis_h2c_tuser_zero_byte; // @[FpgaCloudSerHw.scala 68:26]
  wire  qdma_io_qdma_port_m_axis_h2c_tlast; // @[FpgaCloudSerHw.scala 68:26]
  wire  qdma_io_qdma_port_m_axis_h2c_tvalid; // @[FpgaCloudSerHw.scala 68:26]
  wire  qdma_io_qdma_port_m_axis_h2c_tready; // @[FpgaCloudSerHw.scala 68:26]
  wire  qdma_io_user_clk; // @[FpgaCloudSerHw.scala 68:26]
  wire  qdma_io_user_arstn; // @[FpgaCloudSerHw.scala 68:26]
  wire  qdma_io_h2c_cmd_ready; // @[FpgaCloudSerHw.scala 68:26]
  wire  qdma_io_h2c_cmd_valid; // @[FpgaCloudSerHw.scala 68:26]
  wire [63:0] qdma_io_h2c_cmd_bits_addr; // @[FpgaCloudSerHw.scala 68:26]
  wire [31:0] qdma_io_h2c_cmd_bits_len; // @[FpgaCloudSerHw.scala 68:26]
  wire  qdma_io_h2c_data_valid; // @[FpgaCloudSerHw.scala 68:26]
  wire [31:0] qdma_io_reg_control_0; // @[FpgaCloudSerHw.scala 68:26]
  wire [31:0] qdma_io_reg_control_8; // @[FpgaCloudSerHw.scala 68:26]
  wire [31:0] qdma_io_reg_control_9; // @[FpgaCloudSerHw.scala 68:26]
  wire [31:0] qdma_io_reg_control_10; // @[FpgaCloudSerHw.scala 68:26]
  wire [31:0] qdma_io_reg_control_11; // @[FpgaCloudSerHw.scala 68:26]
  wire [31:0] qdma_io_reg_control_12; // @[FpgaCloudSerHw.scala 68:26]
  wire [31:0] qdma_io_reg_control_13; // @[FpgaCloudSerHw.scala 68:26]
  wire [31:0] qdma_io_reg_control_14; // @[FpgaCloudSerHw.scala 68:26]
  wire [31:0] qdma_io_reg_status_300; // @[FpgaCloudSerHw.scala 68:26]
  wire [31:0] qdma_io_reg_status_400; // @[FpgaCloudSerHw.scala 68:26]
  wire [31:0] qdma_io_reg_status_401; // @[FpgaCloudSerHw.scala 68:26]
  wire [31:0] qdma_io_reg_status_402; // @[FpgaCloudSerHw.scala 68:26]
  wire [31:0] qdma_io_reg_status_403; // @[FpgaCloudSerHw.scala 68:26]
  wire [31:0] qdma_io_reg_status_404; // @[FpgaCloudSerHw.scala 68:26]
  wire [31:0] qdma_io_reg_status_405; // @[FpgaCloudSerHw.scala 68:26]
  wire [31:0] qdma_io_reg_status_406; // @[FpgaCloudSerHw.scala 68:26]
  wire [31:0] qdma_io_reg_status_407; // @[FpgaCloudSerHw.scala 68:26]
  wire [31:0] qdma_io_reg_status_408; // @[FpgaCloudSerHw.scala 68:26]
  wire [31:0] qdma_io_reg_status_409; // @[FpgaCloudSerHw.scala 68:26]
  wire [31:0] qdma_io_reg_status_410; // @[FpgaCloudSerHw.scala 68:26]
  wire [31:0] qdma_io_reg_status_411; // @[FpgaCloudSerHw.scala 68:26]
  wire [31:0] qdma_io_reg_status_412; // @[FpgaCloudSerHw.scala 68:26]
  wire [31:0] qdma_io_reg_status_413; // @[FpgaCloudSerHw.scala 68:26]
  wire [31:0] qdma_io_reg_status_414; // @[FpgaCloudSerHw.scala 68:26]
  wire  qdma_io_axib_aw_ready; // @[FpgaCloudSerHw.scala 68:26]
  wire  qdma_io_axib_aw_valid; // @[FpgaCloudSerHw.scala 68:26]
  wire [63:0] qdma_io_axib_aw_bits_addr; // @[FpgaCloudSerHw.scala 68:26]
  wire  qdma_io_axib_w_ready; // @[FpgaCloudSerHw.scala 68:26]
  wire  qdma_io_axib_w_valid; // @[FpgaCloudSerHw.scala 68:26]
  wire [511:0] qdma_io_axib_w_bits_data; // @[FpgaCloudSerHw.scala 68:26]
  wire  qdma_io_axib_r_ready; // @[FpgaCloudSerHw.scala 68:26]
  wire [511:0] qdma_io_axib_r_bits_data; // @[FpgaCloudSerHw.scala 68:26]
  wire  qdma_io_out_valid; // @[FpgaCloudSerHw.scala 68:26]
  wire [31:0] qdma_counter_4_0; // @[FpgaCloudSerHw.scala 68:26]
  wire  qdma_io_out_ready; // @[FpgaCloudSerHw.scala 68:26]
  wire [31:0] qdma_counter_7_0; // @[FpgaCloudSerHw.scala 68:26]
  wire [31:0] qdma_counter_1_0; // @[FpgaCloudSerHw.scala 68:26]
  wire  qdma_io_in_ready; // @[FpgaCloudSerHw.scala 68:26]
  wire [31:0] qdma_counter_3_1; // @[FpgaCloudSerHw.scala 68:26]
  wire  qdma_io_out_ready_0; // @[FpgaCloudSerHw.scala 68:26]
  wire [31:0] qdma_counter_6_0; // @[FpgaCloudSerHw.scala 68:26]
  wire  qdma_io_out_valid_0; // @[FpgaCloudSerHw.scala 68:26]
  wire [31:0] qdma_counter_0; // @[FpgaCloudSerHw.scala 68:26]
  wire  qdma_io_in_valid; // @[FpgaCloudSerHw.scala 68:26]
  wire [31:0] qdma_io_tlb_miss_count; // @[FpgaCloudSerHw.scala 68:26]
  wire  qdma_io_out_valid_1; // @[FpgaCloudSerHw.scala 68:26]
  wire [31:0] qdma_counter_2_1; // @[FpgaCloudSerHw.scala 68:26]
  wire [31:0] qdma_counter_5_0; // @[FpgaCloudSerHw.scala 68:26]
  wire  qdma_io_out_ready_1; // @[FpgaCloudSerHw.scala 68:26]
  wire  ser_clock; // @[FpgaCloudSerHw.scala 104:21]
  wire  ser_reset; // @[FpgaCloudSerHw.scala 104:21]
  wire  ser_io_meta_in_ready; // @[FpgaCloudSerHw.scala 104:21]
  wire  ser_io_meta_in_valid; // @[FpgaCloudSerHw.scala 104:21]
  wire [9:0] ser_io_meta_in_bits_class_id; // @[FpgaCloudSerHw.scala 104:21]
  wire [63:0] ser_io_meta_in_bits_host_base_addr; // @[FpgaCloudSerHw.scala 104:21]
  wire  ser_io_host_data_in_ready; // @[FpgaCloudSerHw.scala 104:21]
  wire  ser_io_host_data_in_valid; // @[FpgaCloudSerHw.scala 104:21]
  wire  ser_io_host_data_cmd_ready; // @[FpgaCloudSerHw.scala 104:21]
  wire  ser_io_host_data_cmd_valid; // @[FpgaCloudSerHw.scala 104:21]
  wire [63:0] ser_io_host_data_cmd_bits_vaddr; // @[FpgaCloudSerHw.scala 104:21]
  wire [31:0] ser_io_host_data_cmd_bits_length; // @[FpgaCloudSerHw.scala 104:21]
  wire  ser_io_class_meta_req_ready; // @[FpgaCloudSerHw.scala 104:21]
  wire  ser_io_class_meta_req_valid; // @[FpgaCloudSerHw.scala 104:21]
  wire [9:0] ser_io_class_meta_req_bits_class_id; // @[FpgaCloudSerHw.scala 104:21]
  wire  ser_io_class_meta_rsp_valid; // @[FpgaCloudSerHw.scala 104:21]
  wire [7:0] ser_io_class_meta_rsp_bits_class_meta_max_field_num; // @[FpgaCloudSerHw.scala 104:21]
  wire  ser_io_class_meta_rsp_bits_class_meta_field_type_0_is_repeated; // @[FpgaCloudSerHw.scala 104:21]
  wire [4:0] ser_io_class_meta_rsp_bits_class_meta_field_type_0_field_type; // @[FpgaCloudSerHw.scala 104:21]
  wire [15:0] ser_io_class_meta_rsp_bits_class_meta_field_type_0_sub_class_id; // @[FpgaCloudSerHw.scala 104:21]
  wire  ser_io_class_meta_rsp_bits_class_meta_field_type_1_is_repeated; // @[FpgaCloudSerHw.scala 104:21]
  wire [4:0] ser_io_class_meta_rsp_bits_class_meta_field_type_1_field_type; // @[FpgaCloudSerHw.scala 104:21]
  wire [15:0] ser_io_class_meta_rsp_bits_class_meta_field_type_1_sub_class_id; // @[FpgaCloudSerHw.scala 104:21]
  wire  ser_io_class_meta_rsp_bits_class_meta_field_type_2_is_repeated; // @[FpgaCloudSerHw.scala 104:21]
  wire [4:0] ser_io_class_meta_rsp_bits_class_meta_field_type_2_field_type; // @[FpgaCloudSerHw.scala 104:21]
  wire [15:0] ser_io_class_meta_rsp_bits_class_meta_field_type_2_sub_class_id; // @[FpgaCloudSerHw.scala 104:21]
  wire  ser_io_class_meta_rsp_bits_class_meta_field_type_3_is_repeated; // @[FpgaCloudSerHw.scala 104:21]
  wire [4:0] ser_io_class_meta_rsp_bits_class_meta_field_type_3_field_type; // @[FpgaCloudSerHw.scala 104:21]
  wire [15:0] ser_io_class_meta_rsp_bits_class_meta_field_type_3_sub_class_id; // @[FpgaCloudSerHw.scala 104:21]
  wire  ser_io_class_meta_rsp_bits_class_meta_field_type_4_is_repeated; // @[FpgaCloudSerHw.scala 104:21]
  wire [4:0] ser_io_class_meta_rsp_bits_class_meta_field_type_4_field_type; // @[FpgaCloudSerHw.scala 104:21]
  wire [15:0] ser_io_class_meta_rsp_bits_class_meta_field_type_4_sub_class_id; // @[FpgaCloudSerHw.scala 104:21]
  wire  ser_io_class_meta_rsp_bits_class_meta_field_type_5_is_repeated; // @[FpgaCloudSerHw.scala 104:21]
  wire [4:0] ser_io_class_meta_rsp_bits_class_meta_field_type_5_field_type; // @[FpgaCloudSerHw.scala 104:21]
  wire [15:0] ser_io_class_meta_rsp_bits_class_meta_field_type_5_sub_class_id; // @[FpgaCloudSerHw.scala 104:21]
  wire  ser_io_class_meta_rsp_bits_class_meta_field_type_6_is_repeated; // @[FpgaCloudSerHw.scala 104:21]
  wire [4:0] ser_io_class_meta_rsp_bits_class_meta_field_type_6_field_type; // @[FpgaCloudSerHw.scala 104:21]
  wire [15:0] ser_io_class_meta_rsp_bits_class_meta_field_type_6_sub_class_id; // @[FpgaCloudSerHw.scala 104:21]
  wire  ser_io_class_meta_rsp_bits_class_meta_field_type_7_is_repeated; // @[FpgaCloudSerHw.scala 104:21]
  wire [4:0] ser_io_class_meta_rsp_bits_class_meta_field_type_7_field_type; // @[FpgaCloudSerHw.scala 104:21]
  wire [15:0] ser_io_class_meta_rsp_bits_class_meta_field_type_7_sub_class_id; // @[FpgaCloudSerHw.scala 104:21]
  wire  ser_io_class_meta_rsp_bits_class_meta_field_type_8_is_repeated; // @[FpgaCloudSerHw.scala 104:21]
  wire [4:0] ser_io_class_meta_rsp_bits_class_meta_field_type_8_field_type; // @[FpgaCloudSerHw.scala 104:21]
  wire [15:0] ser_io_class_meta_rsp_bits_class_meta_field_type_8_sub_class_id; // @[FpgaCloudSerHw.scala 104:21]
  wire  ser_io_class_meta_rsp_bits_class_meta_field_type_9_is_repeated; // @[FpgaCloudSerHw.scala 104:21]
  wire [4:0] ser_io_class_meta_rsp_bits_class_meta_field_type_9_field_type; // @[FpgaCloudSerHw.scala 104:21]
  wire [15:0] ser_io_class_meta_rsp_bits_class_meta_field_type_9_sub_class_id; // @[FpgaCloudSerHw.scala 104:21]
  wire  ser_io_class_meta_rsp_bits_class_meta_field_type_10_is_repeated; // @[FpgaCloudSerHw.scala 104:21]
  wire [4:0] ser_io_class_meta_rsp_bits_class_meta_field_type_10_field_type; // @[FpgaCloudSerHw.scala 104:21]
  wire [15:0] ser_io_class_meta_rsp_bits_class_meta_field_type_10_sub_class_id; // @[FpgaCloudSerHw.scala 104:21]
  wire  ser_io_class_meta_rsp_bits_class_meta_field_type_11_is_repeated; // @[FpgaCloudSerHw.scala 104:21]
  wire [4:0] ser_io_class_meta_rsp_bits_class_meta_field_type_11_field_type; // @[FpgaCloudSerHw.scala 104:21]
  wire [15:0] ser_io_class_meta_rsp_bits_class_meta_field_type_11_sub_class_id; // @[FpgaCloudSerHw.scala 104:21]
  wire  ser_io_class_meta_rsp_bits_class_meta_field_type_12_is_repeated; // @[FpgaCloudSerHw.scala 104:21]
  wire [4:0] ser_io_class_meta_rsp_bits_class_meta_field_type_12_field_type; // @[FpgaCloudSerHw.scala 104:21]
  wire [15:0] ser_io_class_meta_rsp_bits_class_meta_field_type_12_sub_class_id; // @[FpgaCloudSerHw.scala 104:21]
  wire  ser_io_class_meta_rsp_bits_class_meta_field_type_13_is_repeated; // @[FpgaCloudSerHw.scala 104:21]
  wire [4:0] ser_io_class_meta_rsp_bits_class_meta_field_type_13_field_type; // @[FpgaCloudSerHw.scala 104:21]
  wire [15:0] ser_io_class_meta_rsp_bits_class_meta_field_type_13_sub_class_id; // @[FpgaCloudSerHw.scala 104:21]
  wire  ser_io_class_meta_rsp_bits_class_meta_field_type_14_is_repeated; // @[FpgaCloudSerHw.scala 104:21]
  wire [4:0] ser_io_class_meta_rsp_bits_class_meta_field_type_14_field_type; // @[FpgaCloudSerHw.scala 104:21]
  wire [15:0] ser_io_class_meta_rsp_bits_class_meta_field_type_14_sub_class_id; // @[FpgaCloudSerHw.scala 104:21]
  wire  ser_io_class_meta_rsp_bits_class_meta_field_type_15_is_repeated; // @[FpgaCloudSerHw.scala 104:21]
  wire [4:0] ser_io_class_meta_rsp_bits_class_meta_field_type_15_field_type; // @[FpgaCloudSerHw.scala 104:21]
  wire [15:0] ser_io_class_meta_rsp_bits_class_meta_field_type_15_sub_class_id; // @[FpgaCloudSerHw.scala 104:21]
  wire  ser_io_class_meta_rsp_bits_class_meta_field_type_16_is_repeated; // @[FpgaCloudSerHw.scala 104:21]
  wire [4:0] ser_io_class_meta_rsp_bits_class_meta_field_type_16_field_type; // @[FpgaCloudSerHw.scala 104:21]
  wire [15:0] ser_io_class_meta_rsp_bits_class_meta_field_type_16_sub_class_id; // @[FpgaCloudSerHw.scala 104:21]
  wire  ser_io_class_meta_rsp_bits_class_meta_field_type_17_is_repeated; // @[FpgaCloudSerHw.scala 104:21]
  wire [4:0] ser_io_class_meta_rsp_bits_class_meta_field_type_17_field_type; // @[FpgaCloudSerHw.scala 104:21]
  wire [15:0] ser_io_class_meta_rsp_bits_class_meta_field_type_17_sub_class_id; // @[FpgaCloudSerHw.scala 104:21]
  wire  ser_io_class_meta_rsp_bits_class_meta_field_type_18_is_repeated; // @[FpgaCloudSerHw.scala 104:21]
  wire [4:0] ser_io_class_meta_rsp_bits_class_meta_field_type_18_field_type; // @[FpgaCloudSerHw.scala 104:21]
  wire [15:0] ser_io_class_meta_rsp_bits_class_meta_field_type_18_sub_class_id; // @[FpgaCloudSerHw.scala 104:21]
  wire  ser_io_class_meta_rsp_bits_class_meta_field_type_19_is_repeated; // @[FpgaCloudSerHw.scala 104:21]
  wire [4:0] ser_io_class_meta_rsp_bits_class_meta_field_type_19_field_type; // @[FpgaCloudSerHw.scala 104:21]
  wire [15:0] ser_io_class_meta_rsp_bits_class_meta_field_type_19_sub_class_id; // @[FpgaCloudSerHw.scala 104:21]
  wire  ser_io_class_meta_rsp_bits_class_meta_field_type_20_is_repeated; // @[FpgaCloudSerHw.scala 104:21]
  wire [4:0] ser_io_class_meta_rsp_bits_class_meta_field_type_20_field_type; // @[FpgaCloudSerHw.scala 104:21]
  wire [15:0] ser_io_class_meta_rsp_bits_class_meta_field_type_20_sub_class_id; // @[FpgaCloudSerHw.scala 104:21]
  wire  ser_io_class_meta_rsp_bits_class_meta_field_type_21_is_repeated; // @[FpgaCloudSerHw.scala 104:21]
  wire [4:0] ser_io_class_meta_rsp_bits_class_meta_field_type_21_field_type; // @[FpgaCloudSerHw.scala 104:21]
  wire [15:0] ser_io_class_meta_rsp_bits_class_meta_field_type_21_sub_class_id; // @[FpgaCloudSerHw.scala 104:21]
  wire  ser_io_class_meta_rsp_bits_class_meta_field_type_22_is_repeated; // @[FpgaCloudSerHw.scala 104:21]
  wire [4:0] ser_io_class_meta_rsp_bits_class_meta_field_type_22_field_type; // @[FpgaCloudSerHw.scala 104:21]
  wire [15:0] ser_io_class_meta_rsp_bits_class_meta_field_type_22_sub_class_id; // @[FpgaCloudSerHw.scala 104:21]
  wire  ser_io_class_meta_rsp_bits_class_meta_field_type_23_is_repeated; // @[FpgaCloudSerHw.scala 104:21]
  wire [4:0] ser_io_class_meta_rsp_bits_class_meta_field_type_23_field_type; // @[FpgaCloudSerHw.scala 104:21]
  wire [15:0] ser_io_class_meta_rsp_bits_class_meta_field_type_23_sub_class_id; // @[FpgaCloudSerHw.scala 104:21]
  wire  ser_io_class_meta_rsp_bits_class_meta_field_type_24_is_repeated; // @[FpgaCloudSerHw.scala 104:21]
  wire [4:0] ser_io_class_meta_rsp_bits_class_meta_field_type_24_field_type; // @[FpgaCloudSerHw.scala 104:21]
  wire [15:0] ser_io_class_meta_rsp_bits_class_meta_field_type_24_sub_class_id; // @[FpgaCloudSerHw.scala 104:21]
  wire  ser_io_class_meta_rsp_bits_class_meta_field_type_25_is_repeated; // @[FpgaCloudSerHw.scala 104:21]
  wire [4:0] ser_io_class_meta_rsp_bits_class_meta_field_type_25_field_type; // @[FpgaCloudSerHw.scala 104:21]
  wire [15:0] ser_io_class_meta_rsp_bits_class_meta_field_type_25_sub_class_id; // @[FpgaCloudSerHw.scala 104:21]
  wire  ser_io_class_meta_rsp_bits_class_meta_field_type_26_is_repeated; // @[FpgaCloudSerHw.scala 104:21]
  wire [4:0] ser_io_class_meta_rsp_bits_class_meta_field_type_26_field_type; // @[FpgaCloudSerHw.scala 104:21]
  wire [15:0] ser_io_class_meta_rsp_bits_class_meta_field_type_26_sub_class_id; // @[FpgaCloudSerHw.scala 104:21]
  wire  ser_io_class_meta_rsp_bits_class_meta_field_type_27_is_repeated; // @[FpgaCloudSerHw.scala 104:21]
  wire [4:0] ser_io_class_meta_rsp_bits_class_meta_field_type_27_field_type; // @[FpgaCloudSerHw.scala 104:21]
  wire [15:0] ser_io_class_meta_rsp_bits_class_meta_field_type_27_sub_class_id; // @[FpgaCloudSerHw.scala 104:21]
  wire  ser_io_class_meta_rsp_bits_class_meta_field_type_28_is_repeated; // @[FpgaCloudSerHw.scala 104:21]
  wire [4:0] ser_io_class_meta_rsp_bits_class_meta_field_type_28_field_type; // @[FpgaCloudSerHw.scala 104:21]
  wire [15:0] ser_io_class_meta_rsp_bits_class_meta_field_type_28_sub_class_id; // @[FpgaCloudSerHw.scala 104:21]
  wire  ser_io_class_meta_rsp_bits_class_meta_field_type_29_is_repeated; // @[FpgaCloudSerHw.scala 104:21]
  wire [4:0] ser_io_class_meta_rsp_bits_class_meta_field_type_29_field_type; // @[FpgaCloudSerHw.scala 104:21]
  wire [15:0] ser_io_class_meta_rsp_bits_class_meta_field_type_29_sub_class_id; // @[FpgaCloudSerHw.scala 104:21]
  wire  ser_io_class_meta_rsp_bits_class_meta_field_type_30_is_repeated; // @[FpgaCloudSerHw.scala 104:21]
  wire [4:0] ser_io_class_meta_rsp_bits_class_meta_field_type_30_field_type; // @[FpgaCloudSerHw.scala 104:21]
  wire [15:0] ser_io_class_meta_rsp_bits_class_meta_field_type_30_sub_class_id; // @[FpgaCloudSerHw.scala 104:21]
  wire  ser_io_class_meta_rsp_bits_class_meta_field_type_31_is_repeated; // @[FpgaCloudSerHw.scala 104:21]
  wire [4:0] ser_io_class_meta_rsp_bits_class_meta_field_type_31_field_type; // @[FpgaCloudSerHw.scala 104:21]
  wire [15:0] ser_io_class_meta_rsp_bits_class_meta_field_type_31_sub_class_id; // @[FpgaCloudSerHw.scala 104:21]
  wire  ser_io_class_meta_rsp_bits_class_meta_field_type_32_is_repeated; // @[FpgaCloudSerHw.scala 104:21]
  wire [4:0] ser_io_class_meta_rsp_bits_class_meta_field_type_32_field_type; // @[FpgaCloudSerHw.scala 104:21]
  wire [15:0] ser_io_class_meta_rsp_bits_class_meta_field_type_32_sub_class_id; // @[FpgaCloudSerHw.scala 104:21]
  wire  ser_io_done_ready; // @[FpgaCloudSerHw.scala 104:21]
  wire  ser_io_done_valid; // @[FpgaCloudSerHw.scala 104:21]
  wire [31:0] ser_counter_3_0; // @[FpgaCloudSerHw.scala 104:21]
  wire [31:0] ser_counter_2_0; // @[FpgaCloudSerHw.scala 104:21]
  wire [31:0] ser_counter_8; // @[FpgaCloudSerHw.scala 104:21]
  wire [31:0] ser_counter_1_1; // @[FpgaCloudSerHw.scala 104:21]
  wire  meta_table_clock; // @[FpgaCloudSerHw.scala 105:28]
  wire  meta_table_reset; // @[FpgaCloudSerHw.scala 105:28]
  wire  meta_table_io_class_meta_init_ready; // @[FpgaCloudSerHw.scala 105:28]
  wire  meta_table_io_class_meta_init_valid; // @[FpgaCloudSerHw.scala 105:28]
  wire [9:0] meta_table_io_class_meta_init_bits_class_id; // @[FpgaCloudSerHw.scala 105:28]
  wire [15:0] meta_table_io_class_meta_init_bits_desc_state_class_length; // @[FpgaCloudSerHw.scala 105:28]
  wire [7:0] meta_table_io_class_meta_init_bits_desc_state_max_field_num; // @[FpgaCloudSerHw.scala 105:28]
  wire  meta_table_io_class_meta_init_bits_desc_state_field_type_0_is_repeated; // @[FpgaCloudSerHw.scala 105:28]
  wire [4:0] meta_table_io_class_meta_init_bits_desc_state_field_type_0_field_type; // @[FpgaCloudSerHw.scala 105:28]
  wire [15:0] meta_table_io_class_meta_init_bits_desc_state_field_type_0_sub_class_id; // @[FpgaCloudSerHw.scala 105:28]
  wire  meta_table_io_class_meta_init_bits_desc_state_field_type_0_is_host; // @[FpgaCloudSerHw.scala 105:28]
  wire  meta_table_io_class_meta_init_bits_desc_state_field_type_1_is_repeated; // @[FpgaCloudSerHw.scala 105:28]
  wire [4:0] meta_table_io_class_meta_init_bits_desc_state_field_type_1_field_type; // @[FpgaCloudSerHw.scala 105:28]
  wire [15:0] meta_table_io_class_meta_init_bits_desc_state_field_type_1_sub_class_id; // @[FpgaCloudSerHw.scala 105:28]
  wire  meta_table_io_class_meta_init_bits_desc_state_field_type_1_is_host; // @[FpgaCloudSerHw.scala 105:28]
  wire  meta_table_io_class_meta_init_bits_desc_state_field_type_2_is_repeated; // @[FpgaCloudSerHw.scala 105:28]
  wire [4:0] meta_table_io_class_meta_init_bits_desc_state_field_type_2_field_type; // @[FpgaCloudSerHw.scala 105:28]
  wire [15:0] meta_table_io_class_meta_init_bits_desc_state_field_type_2_sub_class_id; // @[FpgaCloudSerHw.scala 105:28]
  wire  meta_table_io_class_meta_init_bits_desc_state_field_type_2_is_host; // @[FpgaCloudSerHw.scala 105:28]
  wire  meta_table_io_class_meta_init_bits_desc_state_field_type_3_is_repeated; // @[FpgaCloudSerHw.scala 105:28]
  wire [4:0] meta_table_io_class_meta_init_bits_desc_state_field_type_3_field_type; // @[FpgaCloudSerHw.scala 105:28]
  wire [15:0] meta_table_io_class_meta_init_bits_desc_state_field_type_3_sub_class_id; // @[FpgaCloudSerHw.scala 105:28]
  wire  meta_table_io_class_meta_init_bits_desc_state_field_type_3_is_host; // @[FpgaCloudSerHw.scala 105:28]
  wire  meta_table_io_class_meta_init_bits_desc_state_field_type_4_is_repeated; // @[FpgaCloudSerHw.scala 105:28]
  wire [4:0] meta_table_io_class_meta_init_bits_desc_state_field_type_4_field_type; // @[FpgaCloudSerHw.scala 105:28]
  wire [15:0] meta_table_io_class_meta_init_bits_desc_state_field_type_4_sub_class_id; // @[FpgaCloudSerHw.scala 105:28]
  wire  meta_table_io_class_meta_init_bits_desc_state_field_type_4_is_host; // @[FpgaCloudSerHw.scala 105:28]
  wire  meta_table_io_class_meta_init_bits_desc_state_field_type_5_is_repeated; // @[FpgaCloudSerHw.scala 105:28]
  wire [4:0] meta_table_io_class_meta_init_bits_desc_state_field_type_5_field_type; // @[FpgaCloudSerHw.scala 105:28]
  wire [15:0] meta_table_io_class_meta_init_bits_desc_state_field_type_5_sub_class_id; // @[FpgaCloudSerHw.scala 105:28]
  wire  meta_table_io_class_meta_init_bits_desc_state_field_type_5_is_host; // @[FpgaCloudSerHw.scala 105:28]
  wire  meta_table_io_class_meta_init_bits_desc_state_field_type_6_is_repeated; // @[FpgaCloudSerHw.scala 105:28]
  wire [4:0] meta_table_io_class_meta_init_bits_desc_state_field_type_6_field_type; // @[FpgaCloudSerHw.scala 105:28]
  wire [15:0] meta_table_io_class_meta_init_bits_desc_state_field_type_6_sub_class_id; // @[FpgaCloudSerHw.scala 105:28]
  wire  meta_table_io_class_meta_init_bits_desc_state_field_type_6_is_host; // @[FpgaCloudSerHw.scala 105:28]
  wire  meta_table_io_class_meta_init_bits_desc_state_field_type_7_is_repeated; // @[FpgaCloudSerHw.scala 105:28]
  wire [4:0] meta_table_io_class_meta_init_bits_desc_state_field_type_7_field_type; // @[FpgaCloudSerHw.scala 105:28]
  wire [15:0] meta_table_io_class_meta_init_bits_desc_state_field_type_7_sub_class_id; // @[FpgaCloudSerHw.scala 105:28]
  wire  meta_table_io_class_meta_init_bits_desc_state_field_type_7_is_host; // @[FpgaCloudSerHw.scala 105:28]
  wire  meta_table_io_class_meta_init_bits_desc_state_field_type_8_is_repeated; // @[FpgaCloudSerHw.scala 105:28]
  wire [4:0] meta_table_io_class_meta_init_bits_desc_state_field_type_8_field_type; // @[FpgaCloudSerHw.scala 105:28]
  wire [15:0] meta_table_io_class_meta_init_bits_desc_state_field_type_8_sub_class_id; // @[FpgaCloudSerHw.scala 105:28]
  wire  meta_table_io_class_meta_init_bits_desc_state_field_type_8_is_host; // @[FpgaCloudSerHw.scala 105:28]
  wire  meta_table_io_class_meta_init_bits_desc_state_field_type_9_is_repeated; // @[FpgaCloudSerHw.scala 105:28]
  wire [4:0] meta_table_io_class_meta_init_bits_desc_state_field_type_9_field_type; // @[FpgaCloudSerHw.scala 105:28]
  wire [15:0] meta_table_io_class_meta_init_bits_desc_state_field_type_9_sub_class_id; // @[FpgaCloudSerHw.scala 105:28]
  wire  meta_table_io_class_meta_init_bits_desc_state_field_type_9_is_host; // @[FpgaCloudSerHw.scala 105:28]
  wire  meta_table_io_class_meta_init_bits_desc_state_field_type_10_is_repeated; // @[FpgaCloudSerHw.scala 105:28]
  wire [4:0] meta_table_io_class_meta_init_bits_desc_state_field_type_10_field_type; // @[FpgaCloudSerHw.scala 105:28]
  wire [15:0] meta_table_io_class_meta_init_bits_desc_state_field_type_10_sub_class_id; // @[FpgaCloudSerHw.scala 105:28]
  wire  meta_table_io_class_meta_init_bits_desc_state_field_type_10_is_host; // @[FpgaCloudSerHw.scala 105:28]
  wire  meta_table_io_class_meta_init_bits_desc_state_field_type_11_is_repeated; // @[FpgaCloudSerHw.scala 105:28]
  wire [4:0] meta_table_io_class_meta_init_bits_desc_state_field_type_11_field_type; // @[FpgaCloudSerHw.scala 105:28]
  wire [15:0] meta_table_io_class_meta_init_bits_desc_state_field_type_11_sub_class_id; // @[FpgaCloudSerHw.scala 105:28]
  wire  meta_table_io_class_meta_init_bits_desc_state_field_type_11_is_host; // @[FpgaCloudSerHw.scala 105:28]
  wire  meta_table_io_class_meta_init_bits_desc_state_field_type_12_is_repeated; // @[FpgaCloudSerHw.scala 105:28]
  wire [4:0] meta_table_io_class_meta_init_bits_desc_state_field_type_12_field_type; // @[FpgaCloudSerHw.scala 105:28]
  wire [15:0] meta_table_io_class_meta_init_bits_desc_state_field_type_12_sub_class_id; // @[FpgaCloudSerHw.scala 105:28]
  wire  meta_table_io_class_meta_init_bits_desc_state_field_type_12_is_host; // @[FpgaCloudSerHw.scala 105:28]
  wire  meta_table_io_class_meta_init_bits_desc_state_field_type_13_is_repeated; // @[FpgaCloudSerHw.scala 105:28]
  wire [4:0] meta_table_io_class_meta_init_bits_desc_state_field_type_13_field_type; // @[FpgaCloudSerHw.scala 105:28]
  wire [15:0] meta_table_io_class_meta_init_bits_desc_state_field_type_13_sub_class_id; // @[FpgaCloudSerHw.scala 105:28]
  wire  meta_table_io_class_meta_init_bits_desc_state_field_type_13_is_host; // @[FpgaCloudSerHw.scala 105:28]
  wire  meta_table_io_class_meta_init_bits_desc_state_field_type_14_is_repeated; // @[FpgaCloudSerHw.scala 105:28]
  wire [4:0] meta_table_io_class_meta_init_bits_desc_state_field_type_14_field_type; // @[FpgaCloudSerHw.scala 105:28]
  wire [15:0] meta_table_io_class_meta_init_bits_desc_state_field_type_14_sub_class_id; // @[FpgaCloudSerHw.scala 105:28]
  wire  meta_table_io_class_meta_init_bits_desc_state_field_type_14_is_host; // @[FpgaCloudSerHw.scala 105:28]
  wire  meta_table_io_class_meta_init_bits_desc_state_field_type_15_is_repeated; // @[FpgaCloudSerHw.scala 105:28]
  wire [4:0] meta_table_io_class_meta_init_bits_desc_state_field_type_15_field_type; // @[FpgaCloudSerHw.scala 105:28]
  wire [15:0] meta_table_io_class_meta_init_bits_desc_state_field_type_15_sub_class_id; // @[FpgaCloudSerHw.scala 105:28]
  wire  meta_table_io_class_meta_init_bits_desc_state_field_type_15_is_host; // @[FpgaCloudSerHw.scala 105:28]
  wire  meta_table_io_class_meta_init_bits_desc_state_field_type_16_is_repeated; // @[FpgaCloudSerHw.scala 105:28]
  wire [4:0] meta_table_io_class_meta_init_bits_desc_state_field_type_16_field_type; // @[FpgaCloudSerHw.scala 105:28]
  wire [15:0] meta_table_io_class_meta_init_bits_desc_state_field_type_16_sub_class_id; // @[FpgaCloudSerHw.scala 105:28]
  wire  meta_table_io_class_meta_init_bits_desc_state_field_type_16_is_host; // @[FpgaCloudSerHw.scala 105:28]
  wire  meta_table_io_class_meta_init_bits_desc_state_field_type_17_is_repeated; // @[FpgaCloudSerHw.scala 105:28]
  wire [4:0] meta_table_io_class_meta_init_bits_desc_state_field_type_17_field_type; // @[FpgaCloudSerHw.scala 105:28]
  wire [15:0] meta_table_io_class_meta_init_bits_desc_state_field_type_17_sub_class_id; // @[FpgaCloudSerHw.scala 105:28]
  wire  meta_table_io_class_meta_init_bits_desc_state_field_type_17_is_host; // @[FpgaCloudSerHw.scala 105:28]
  wire  meta_table_io_class_meta_init_bits_desc_state_field_type_18_is_repeated; // @[FpgaCloudSerHw.scala 105:28]
  wire [4:0] meta_table_io_class_meta_init_bits_desc_state_field_type_18_field_type; // @[FpgaCloudSerHw.scala 105:28]
  wire [15:0] meta_table_io_class_meta_init_bits_desc_state_field_type_18_sub_class_id; // @[FpgaCloudSerHw.scala 105:28]
  wire  meta_table_io_class_meta_init_bits_desc_state_field_type_18_is_host; // @[FpgaCloudSerHw.scala 105:28]
  wire  meta_table_io_class_meta_init_bits_desc_state_field_type_19_is_repeated; // @[FpgaCloudSerHw.scala 105:28]
  wire [4:0] meta_table_io_class_meta_init_bits_desc_state_field_type_19_field_type; // @[FpgaCloudSerHw.scala 105:28]
  wire [15:0] meta_table_io_class_meta_init_bits_desc_state_field_type_19_sub_class_id; // @[FpgaCloudSerHw.scala 105:28]
  wire  meta_table_io_class_meta_init_bits_desc_state_field_type_19_is_host; // @[FpgaCloudSerHw.scala 105:28]
  wire  meta_table_io_class_meta_init_bits_desc_state_field_type_20_is_repeated; // @[FpgaCloudSerHw.scala 105:28]
  wire [4:0] meta_table_io_class_meta_init_bits_desc_state_field_type_20_field_type; // @[FpgaCloudSerHw.scala 105:28]
  wire [15:0] meta_table_io_class_meta_init_bits_desc_state_field_type_20_sub_class_id; // @[FpgaCloudSerHw.scala 105:28]
  wire  meta_table_io_class_meta_init_bits_desc_state_field_type_20_is_host; // @[FpgaCloudSerHw.scala 105:28]
  wire  meta_table_io_class_meta_init_bits_desc_state_field_type_21_is_repeated; // @[FpgaCloudSerHw.scala 105:28]
  wire [4:0] meta_table_io_class_meta_init_bits_desc_state_field_type_21_field_type; // @[FpgaCloudSerHw.scala 105:28]
  wire [15:0] meta_table_io_class_meta_init_bits_desc_state_field_type_21_sub_class_id; // @[FpgaCloudSerHw.scala 105:28]
  wire  meta_table_io_class_meta_init_bits_desc_state_field_type_21_is_host; // @[FpgaCloudSerHw.scala 105:28]
  wire  meta_table_io_class_meta_init_bits_desc_state_field_type_22_is_repeated; // @[FpgaCloudSerHw.scala 105:28]
  wire [4:0] meta_table_io_class_meta_init_bits_desc_state_field_type_22_field_type; // @[FpgaCloudSerHw.scala 105:28]
  wire [15:0] meta_table_io_class_meta_init_bits_desc_state_field_type_22_sub_class_id; // @[FpgaCloudSerHw.scala 105:28]
  wire  meta_table_io_class_meta_init_bits_desc_state_field_type_22_is_host; // @[FpgaCloudSerHw.scala 105:28]
  wire  meta_table_io_class_meta_init_bits_desc_state_field_type_23_is_repeated; // @[FpgaCloudSerHw.scala 105:28]
  wire [4:0] meta_table_io_class_meta_init_bits_desc_state_field_type_23_field_type; // @[FpgaCloudSerHw.scala 105:28]
  wire [15:0] meta_table_io_class_meta_init_bits_desc_state_field_type_23_sub_class_id; // @[FpgaCloudSerHw.scala 105:28]
  wire  meta_table_io_class_meta_init_bits_desc_state_field_type_23_is_host; // @[FpgaCloudSerHw.scala 105:28]
  wire  meta_table_io_class_meta_init_bits_desc_state_field_type_24_is_repeated; // @[FpgaCloudSerHw.scala 105:28]
  wire [4:0] meta_table_io_class_meta_init_bits_desc_state_field_type_24_field_type; // @[FpgaCloudSerHw.scala 105:28]
  wire [15:0] meta_table_io_class_meta_init_bits_desc_state_field_type_24_sub_class_id; // @[FpgaCloudSerHw.scala 105:28]
  wire  meta_table_io_class_meta_init_bits_desc_state_field_type_24_is_host; // @[FpgaCloudSerHw.scala 105:28]
  wire  meta_table_io_class_meta_init_bits_desc_state_field_type_25_is_repeated; // @[FpgaCloudSerHw.scala 105:28]
  wire [4:0] meta_table_io_class_meta_init_bits_desc_state_field_type_25_field_type; // @[FpgaCloudSerHw.scala 105:28]
  wire [15:0] meta_table_io_class_meta_init_bits_desc_state_field_type_25_sub_class_id; // @[FpgaCloudSerHw.scala 105:28]
  wire  meta_table_io_class_meta_init_bits_desc_state_field_type_25_is_host; // @[FpgaCloudSerHw.scala 105:28]
  wire  meta_table_io_class_meta_init_bits_desc_state_field_type_26_is_repeated; // @[FpgaCloudSerHw.scala 105:28]
  wire [4:0] meta_table_io_class_meta_init_bits_desc_state_field_type_26_field_type; // @[FpgaCloudSerHw.scala 105:28]
  wire [15:0] meta_table_io_class_meta_init_bits_desc_state_field_type_26_sub_class_id; // @[FpgaCloudSerHw.scala 105:28]
  wire  meta_table_io_class_meta_init_bits_desc_state_field_type_26_is_host; // @[FpgaCloudSerHw.scala 105:28]
  wire  meta_table_io_class_meta_init_bits_desc_state_field_type_27_is_repeated; // @[FpgaCloudSerHw.scala 105:28]
  wire [4:0] meta_table_io_class_meta_init_bits_desc_state_field_type_27_field_type; // @[FpgaCloudSerHw.scala 105:28]
  wire [15:0] meta_table_io_class_meta_init_bits_desc_state_field_type_27_sub_class_id; // @[FpgaCloudSerHw.scala 105:28]
  wire  meta_table_io_class_meta_init_bits_desc_state_field_type_27_is_host; // @[FpgaCloudSerHw.scala 105:28]
  wire  meta_table_io_class_meta_init_bits_desc_state_field_type_28_is_repeated; // @[FpgaCloudSerHw.scala 105:28]
  wire [4:0] meta_table_io_class_meta_init_bits_desc_state_field_type_28_field_type; // @[FpgaCloudSerHw.scala 105:28]
  wire [15:0] meta_table_io_class_meta_init_bits_desc_state_field_type_28_sub_class_id; // @[FpgaCloudSerHw.scala 105:28]
  wire  meta_table_io_class_meta_init_bits_desc_state_field_type_28_is_host; // @[FpgaCloudSerHw.scala 105:28]
  wire  meta_table_io_class_meta_init_bits_desc_state_field_type_29_is_repeated; // @[FpgaCloudSerHw.scala 105:28]
  wire [4:0] meta_table_io_class_meta_init_bits_desc_state_field_type_29_field_type; // @[FpgaCloudSerHw.scala 105:28]
  wire [15:0] meta_table_io_class_meta_init_bits_desc_state_field_type_29_sub_class_id; // @[FpgaCloudSerHw.scala 105:28]
  wire  meta_table_io_class_meta_init_bits_desc_state_field_type_29_is_host; // @[FpgaCloudSerHw.scala 105:28]
  wire  meta_table_io_class_meta_init_bits_desc_state_field_type_30_is_repeated; // @[FpgaCloudSerHw.scala 105:28]
  wire [4:0] meta_table_io_class_meta_init_bits_desc_state_field_type_30_field_type; // @[FpgaCloudSerHw.scala 105:28]
  wire [15:0] meta_table_io_class_meta_init_bits_desc_state_field_type_30_sub_class_id; // @[FpgaCloudSerHw.scala 105:28]
  wire  meta_table_io_class_meta_init_bits_desc_state_field_type_30_is_host; // @[FpgaCloudSerHw.scala 105:28]
  wire  meta_table_io_class_meta_init_bits_desc_state_field_type_31_is_repeated; // @[FpgaCloudSerHw.scala 105:28]
  wire [4:0] meta_table_io_class_meta_init_bits_desc_state_field_type_31_field_type; // @[FpgaCloudSerHw.scala 105:28]
  wire [15:0] meta_table_io_class_meta_init_bits_desc_state_field_type_31_sub_class_id; // @[FpgaCloudSerHw.scala 105:28]
  wire  meta_table_io_class_meta_init_bits_desc_state_field_type_31_is_host; // @[FpgaCloudSerHw.scala 105:28]
  wire  meta_table_io_class_meta_init_bits_desc_state_field_type_32_is_repeated; // @[FpgaCloudSerHw.scala 105:28]
  wire [4:0] meta_table_io_class_meta_init_bits_desc_state_field_type_32_field_type; // @[FpgaCloudSerHw.scala 105:28]
  wire [15:0] meta_table_io_class_meta_init_bits_desc_state_field_type_32_sub_class_id; // @[FpgaCloudSerHw.scala 105:28]
  wire  meta_table_io_class_meta_init_bits_desc_state_field_type_32_is_host; // @[FpgaCloudSerHw.scala 105:28]
  wire  meta_table_io_s_class_meta_req_ready; // @[FpgaCloudSerHw.scala 105:28]
  wire  meta_table_io_s_class_meta_req_valid; // @[FpgaCloudSerHw.scala 105:28]
  wire [9:0] meta_table_io_s_class_meta_req_bits_class_id; // @[FpgaCloudSerHw.scala 105:28]
  wire  meta_table_io_s_class_meta_rsp_valid; // @[FpgaCloudSerHw.scala 105:28]
  wire [7:0] meta_table_io_s_class_meta_rsp_bits_class_meta_max_field_num; // @[FpgaCloudSerHw.scala 105:28]
  wire  meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_0_is_repeated; // @[FpgaCloudSerHw.scala 105:28]
  wire [4:0] meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_0_field_type; // @[FpgaCloudSerHw.scala 105:28]
  wire [15:0] meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_0_sub_class_id; // @[FpgaCloudSerHw.scala 105:28]
  wire  meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_1_is_repeated; // @[FpgaCloudSerHw.scala 105:28]
  wire [4:0] meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_1_field_type; // @[FpgaCloudSerHw.scala 105:28]
  wire [15:0] meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_1_sub_class_id; // @[FpgaCloudSerHw.scala 105:28]
  wire  meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_2_is_repeated; // @[FpgaCloudSerHw.scala 105:28]
  wire [4:0] meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_2_field_type; // @[FpgaCloudSerHw.scala 105:28]
  wire [15:0] meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_2_sub_class_id; // @[FpgaCloudSerHw.scala 105:28]
  wire  meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_3_is_repeated; // @[FpgaCloudSerHw.scala 105:28]
  wire [4:0] meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_3_field_type; // @[FpgaCloudSerHw.scala 105:28]
  wire [15:0] meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_3_sub_class_id; // @[FpgaCloudSerHw.scala 105:28]
  wire  meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_4_is_repeated; // @[FpgaCloudSerHw.scala 105:28]
  wire [4:0] meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_4_field_type; // @[FpgaCloudSerHw.scala 105:28]
  wire [15:0] meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_4_sub_class_id; // @[FpgaCloudSerHw.scala 105:28]
  wire  meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_5_is_repeated; // @[FpgaCloudSerHw.scala 105:28]
  wire [4:0] meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_5_field_type; // @[FpgaCloudSerHw.scala 105:28]
  wire [15:0] meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_5_sub_class_id; // @[FpgaCloudSerHw.scala 105:28]
  wire  meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_6_is_repeated; // @[FpgaCloudSerHw.scala 105:28]
  wire [4:0] meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_6_field_type; // @[FpgaCloudSerHw.scala 105:28]
  wire [15:0] meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_6_sub_class_id; // @[FpgaCloudSerHw.scala 105:28]
  wire  meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_7_is_repeated; // @[FpgaCloudSerHw.scala 105:28]
  wire [4:0] meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_7_field_type; // @[FpgaCloudSerHw.scala 105:28]
  wire [15:0] meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_7_sub_class_id; // @[FpgaCloudSerHw.scala 105:28]
  wire  meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_8_is_repeated; // @[FpgaCloudSerHw.scala 105:28]
  wire [4:0] meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_8_field_type; // @[FpgaCloudSerHw.scala 105:28]
  wire [15:0] meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_8_sub_class_id; // @[FpgaCloudSerHw.scala 105:28]
  wire  meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_9_is_repeated; // @[FpgaCloudSerHw.scala 105:28]
  wire [4:0] meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_9_field_type; // @[FpgaCloudSerHw.scala 105:28]
  wire [15:0] meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_9_sub_class_id; // @[FpgaCloudSerHw.scala 105:28]
  wire  meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_10_is_repeated; // @[FpgaCloudSerHw.scala 105:28]
  wire [4:0] meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_10_field_type; // @[FpgaCloudSerHw.scala 105:28]
  wire [15:0] meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_10_sub_class_id; // @[FpgaCloudSerHw.scala 105:28]
  wire  meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_11_is_repeated; // @[FpgaCloudSerHw.scala 105:28]
  wire [4:0] meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_11_field_type; // @[FpgaCloudSerHw.scala 105:28]
  wire [15:0] meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_11_sub_class_id; // @[FpgaCloudSerHw.scala 105:28]
  wire  meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_12_is_repeated; // @[FpgaCloudSerHw.scala 105:28]
  wire [4:0] meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_12_field_type; // @[FpgaCloudSerHw.scala 105:28]
  wire [15:0] meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_12_sub_class_id; // @[FpgaCloudSerHw.scala 105:28]
  wire  meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_13_is_repeated; // @[FpgaCloudSerHw.scala 105:28]
  wire [4:0] meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_13_field_type; // @[FpgaCloudSerHw.scala 105:28]
  wire [15:0] meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_13_sub_class_id; // @[FpgaCloudSerHw.scala 105:28]
  wire  meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_14_is_repeated; // @[FpgaCloudSerHw.scala 105:28]
  wire [4:0] meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_14_field_type; // @[FpgaCloudSerHw.scala 105:28]
  wire [15:0] meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_14_sub_class_id; // @[FpgaCloudSerHw.scala 105:28]
  wire  meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_15_is_repeated; // @[FpgaCloudSerHw.scala 105:28]
  wire [4:0] meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_15_field_type; // @[FpgaCloudSerHw.scala 105:28]
  wire [15:0] meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_15_sub_class_id; // @[FpgaCloudSerHw.scala 105:28]
  wire  meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_16_is_repeated; // @[FpgaCloudSerHw.scala 105:28]
  wire [4:0] meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_16_field_type; // @[FpgaCloudSerHw.scala 105:28]
  wire [15:0] meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_16_sub_class_id; // @[FpgaCloudSerHw.scala 105:28]
  wire  meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_17_is_repeated; // @[FpgaCloudSerHw.scala 105:28]
  wire [4:0] meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_17_field_type; // @[FpgaCloudSerHw.scala 105:28]
  wire [15:0] meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_17_sub_class_id; // @[FpgaCloudSerHw.scala 105:28]
  wire  meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_18_is_repeated; // @[FpgaCloudSerHw.scala 105:28]
  wire [4:0] meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_18_field_type; // @[FpgaCloudSerHw.scala 105:28]
  wire [15:0] meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_18_sub_class_id; // @[FpgaCloudSerHw.scala 105:28]
  wire  meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_19_is_repeated; // @[FpgaCloudSerHw.scala 105:28]
  wire [4:0] meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_19_field_type; // @[FpgaCloudSerHw.scala 105:28]
  wire [15:0] meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_19_sub_class_id; // @[FpgaCloudSerHw.scala 105:28]
  wire  meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_20_is_repeated; // @[FpgaCloudSerHw.scala 105:28]
  wire [4:0] meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_20_field_type; // @[FpgaCloudSerHw.scala 105:28]
  wire [15:0] meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_20_sub_class_id; // @[FpgaCloudSerHw.scala 105:28]
  wire  meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_21_is_repeated; // @[FpgaCloudSerHw.scala 105:28]
  wire [4:0] meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_21_field_type; // @[FpgaCloudSerHw.scala 105:28]
  wire [15:0] meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_21_sub_class_id; // @[FpgaCloudSerHw.scala 105:28]
  wire  meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_22_is_repeated; // @[FpgaCloudSerHw.scala 105:28]
  wire [4:0] meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_22_field_type; // @[FpgaCloudSerHw.scala 105:28]
  wire [15:0] meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_22_sub_class_id; // @[FpgaCloudSerHw.scala 105:28]
  wire  meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_23_is_repeated; // @[FpgaCloudSerHw.scala 105:28]
  wire [4:0] meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_23_field_type; // @[FpgaCloudSerHw.scala 105:28]
  wire [15:0] meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_23_sub_class_id; // @[FpgaCloudSerHw.scala 105:28]
  wire  meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_24_is_repeated; // @[FpgaCloudSerHw.scala 105:28]
  wire [4:0] meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_24_field_type; // @[FpgaCloudSerHw.scala 105:28]
  wire [15:0] meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_24_sub_class_id; // @[FpgaCloudSerHw.scala 105:28]
  wire  meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_25_is_repeated; // @[FpgaCloudSerHw.scala 105:28]
  wire [4:0] meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_25_field_type; // @[FpgaCloudSerHw.scala 105:28]
  wire [15:0] meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_25_sub_class_id; // @[FpgaCloudSerHw.scala 105:28]
  wire  meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_26_is_repeated; // @[FpgaCloudSerHw.scala 105:28]
  wire [4:0] meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_26_field_type; // @[FpgaCloudSerHw.scala 105:28]
  wire [15:0] meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_26_sub_class_id; // @[FpgaCloudSerHw.scala 105:28]
  wire  meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_27_is_repeated; // @[FpgaCloudSerHw.scala 105:28]
  wire [4:0] meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_27_field_type; // @[FpgaCloudSerHw.scala 105:28]
  wire [15:0] meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_27_sub_class_id; // @[FpgaCloudSerHw.scala 105:28]
  wire  meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_28_is_repeated; // @[FpgaCloudSerHw.scala 105:28]
  wire [4:0] meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_28_field_type; // @[FpgaCloudSerHw.scala 105:28]
  wire [15:0] meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_28_sub_class_id; // @[FpgaCloudSerHw.scala 105:28]
  wire  meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_29_is_repeated; // @[FpgaCloudSerHw.scala 105:28]
  wire [4:0] meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_29_field_type; // @[FpgaCloudSerHw.scala 105:28]
  wire [15:0] meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_29_sub_class_id; // @[FpgaCloudSerHw.scala 105:28]
  wire  meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_30_is_repeated; // @[FpgaCloudSerHw.scala 105:28]
  wire [4:0] meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_30_field_type; // @[FpgaCloudSerHw.scala 105:28]
  wire [15:0] meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_30_sub_class_id; // @[FpgaCloudSerHw.scala 105:28]
  wire  meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_31_is_repeated; // @[FpgaCloudSerHw.scala 105:28]
  wire [4:0] meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_31_field_type; // @[FpgaCloudSerHw.scala 105:28]
  wire [15:0] meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_31_sub_class_id; // @[FpgaCloudSerHw.scala 105:28]
  wire  meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_32_is_repeated; // @[FpgaCloudSerHw.scala 105:28]
  wire [4:0] meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_32_field_type; // @[FpgaCloudSerHw.scala 105:28]
  wire [15:0] meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_32_sub_class_id; // @[FpgaCloudSerHw.scala 105:28]
  wire [31:0] meta_table_counter_5; // @[FpgaCloudSerHw.scala 105:28]
  wire  control_clock; // @[FpgaCloudSerHw.scala 108:29]
  wire  control_reset; // @[FpgaCloudSerHw.scala 108:29]
  wire  control_io_axi_aw_ready; // @[FpgaCloudSerHw.scala 108:29]
  wire  control_io_axi_aw_valid; // @[FpgaCloudSerHw.scala 108:29]
  wire [63:0] control_io_axi_aw_bits_addr; // @[FpgaCloudSerHw.scala 108:29]
  wire  control_io_axi_w_ready; // @[FpgaCloudSerHw.scala 108:29]
  wire  control_io_axi_w_valid; // @[FpgaCloudSerHw.scala 108:29]
  wire [511:0] control_io_axi_w_bits_data; // @[FpgaCloudSerHw.scala 108:29]
  wire  control_io_axi_r_ready; // @[FpgaCloudSerHw.scala 108:29]
  wire  control_io_axi_r_valid; // @[FpgaCloudSerHw.scala 108:29]
  wire [511:0] control_io_axi_r_bits_data; // @[FpgaCloudSerHw.scala 108:29]
  wire  control_io_metadata_init_valid; // @[FpgaCloudSerHw.scala 108:29]
  wire [9:0] control_io_metadata_init_bits_class_id; // @[FpgaCloudSerHw.scala 108:29]
  wire [15:0] control_io_metadata_init_bits_desc_state_class_length; // @[FpgaCloudSerHw.scala 108:29]
  wire [7:0] control_io_metadata_init_bits_desc_state_max_field_num; // @[FpgaCloudSerHw.scala 108:29]
  wire  control_io_metadata_init_bits_desc_state_field_type_0_is_repeated; // @[FpgaCloudSerHw.scala 108:29]
  wire [4:0] control_io_metadata_init_bits_desc_state_field_type_0_field_type; // @[FpgaCloudSerHw.scala 108:29]
  wire [15:0] control_io_metadata_init_bits_desc_state_field_type_0_sub_class_id; // @[FpgaCloudSerHw.scala 108:29]
  wire  control_io_metadata_init_bits_desc_state_field_type_0_is_host; // @[FpgaCloudSerHw.scala 108:29]
  wire  control_io_metadata_init_bits_desc_state_field_type_1_is_repeated; // @[FpgaCloudSerHw.scala 108:29]
  wire [4:0] control_io_metadata_init_bits_desc_state_field_type_1_field_type; // @[FpgaCloudSerHw.scala 108:29]
  wire [15:0] control_io_metadata_init_bits_desc_state_field_type_1_sub_class_id; // @[FpgaCloudSerHw.scala 108:29]
  wire  control_io_metadata_init_bits_desc_state_field_type_1_is_host; // @[FpgaCloudSerHw.scala 108:29]
  wire  control_io_metadata_init_bits_desc_state_field_type_2_is_repeated; // @[FpgaCloudSerHw.scala 108:29]
  wire [4:0] control_io_metadata_init_bits_desc_state_field_type_2_field_type; // @[FpgaCloudSerHw.scala 108:29]
  wire [15:0] control_io_metadata_init_bits_desc_state_field_type_2_sub_class_id; // @[FpgaCloudSerHw.scala 108:29]
  wire  control_io_metadata_init_bits_desc_state_field_type_2_is_host; // @[FpgaCloudSerHw.scala 108:29]
  wire  control_io_metadata_init_bits_desc_state_field_type_3_is_repeated; // @[FpgaCloudSerHw.scala 108:29]
  wire [4:0] control_io_metadata_init_bits_desc_state_field_type_3_field_type; // @[FpgaCloudSerHw.scala 108:29]
  wire [15:0] control_io_metadata_init_bits_desc_state_field_type_3_sub_class_id; // @[FpgaCloudSerHw.scala 108:29]
  wire  control_io_metadata_init_bits_desc_state_field_type_3_is_host; // @[FpgaCloudSerHw.scala 108:29]
  wire  control_io_metadata_init_bits_desc_state_field_type_4_is_repeated; // @[FpgaCloudSerHw.scala 108:29]
  wire [4:0] control_io_metadata_init_bits_desc_state_field_type_4_field_type; // @[FpgaCloudSerHw.scala 108:29]
  wire [15:0] control_io_metadata_init_bits_desc_state_field_type_4_sub_class_id; // @[FpgaCloudSerHw.scala 108:29]
  wire  control_io_metadata_init_bits_desc_state_field_type_4_is_host; // @[FpgaCloudSerHw.scala 108:29]
  wire  control_io_metadata_init_bits_desc_state_field_type_5_is_repeated; // @[FpgaCloudSerHw.scala 108:29]
  wire [4:0] control_io_metadata_init_bits_desc_state_field_type_5_field_type; // @[FpgaCloudSerHw.scala 108:29]
  wire [15:0] control_io_metadata_init_bits_desc_state_field_type_5_sub_class_id; // @[FpgaCloudSerHw.scala 108:29]
  wire  control_io_metadata_init_bits_desc_state_field_type_5_is_host; // @[FpgaCloudSerHw.scala 108:29]
  wire  control_io_metadata_init_bits_desc_state_field_type_6_is_repeated; // @[FpgaCloudSerHw.scala 108:29]
  wire [4:0] control_io_metadata_init_bits_desc_state_field_type_6_field_type; // @[FpgaCloudSerHw.scala 108:29]
  wire [15:0] control_io_metadata_init_bits_desc_state_field_type_6_sub_class_id; // @[FpgaCloudSerHw.scala 108:29]
  wire  control_io_metadata_init_bits_desc_state_field_type_6_is_host; // @[FpgaCloudSerHw.scala 108:29]
  wire  control_io_metadata_init_bits_desc_state_field_type_7_is_repeated; // @[FpgaCloudSerHw.scala 108:29]
  wire [4:0] control_io_metadata_init_bits_desc_state_field_type_7_field_type; // @[FpgaCloudSerHw.scala 108:29]
  wire [15:0] control_io_metadata_init_bits_desc_state_field_type_7_sub_class_id; // @[FpgaCloudSerHw.scala 108:29]
  wire  control_io_metadata_init_bits_desc_state_field_type_7_is_host; // @[FpgaCloudSerHw.scala 108:29]
  wire  control_io_metadata_init_bits_desc_state_field_type_8_is_repeated; // @[FpgaCloudSerHw.scala 108:29]
  wire [4:0] control_io_metadata_init_bits_desc_state_field_type_8_field_type; // @[FpgaCloudSerHw.scala 108:29]
  wire [15:0] control_io_metadata_init_bits_desc_state_field_type_8_sub_class_id; // @[FpgaCloudSerHw.scala 108:29]
  wire  control_io_metadata_init_bits_desc_state_field_type_8_is_host; // @[FpgaCloudSerHw.scala 108:29]
  wire  control_io_metadata_init_bits_desc_state_field_type_9_is_repeated; // @[FpgaCloudSerHw.scala 108:29]
  wire [4:0] control_io_metadata_init_bits_desc_state_field_type_9_field_type; // @[FpgaCloudSerHw.scala 108:29]
  wire [15:0] control_io_metadata_init_bits_desc_state_field_type_9_sub_class_id; // @[FpgaCloudSerHw.scala 108:29]
  wire  control_io_metadata_init_bits_desc_state_field_type_9_is_host; // @[FpgaCloudSerHw.scala 108:29]
  wire  control_io_metadata_init_bits_desc_state_field_type_10_is_repeated; // @[FpgaCloudSerHw.scala 108:29]
  wire [4:0] control_io_metadata_init_bits_desc_state_field_type_10_field_type; // @[FpgaCloudSerHw.scala 108:29]
  wire [15:0] control_io_metadata_init_bits_desc_state_field_type_10_sub_class_id; // @[FpgaCloudSerHw.scala 108:29]
  wire  control_io_metadata_init_bits_desc_state_field_type_10_is_host; // @[FpgaCloudSerHw.scala 108:29]
  wire  control_io_metadata_init_bits_desc_state_field_type_11_is_repeated; // @[FpgaCloudSerHw.scala 108:29]
  wire [4:0] control_io_metadata_init_bits_desc_state_field_type_11_field_type; // @[FpgaCloudSerHw.scala 108:29]
  wire [15:0] control_io_metadata_init_bits_desc_state_field_type_11_sub_class_id; // @[FpgaCloudSerHw.scala 108:29]
  wire  control_io_metadata_init_bits_desc_state_field_type_11_is_host; // @[FpgaCloudSerHw.scala 108:29]
  wire  control_io_metadata_init_bits_desc_state_field_type_12_is_repeated; // @[FpgaCloudSerHw.scala 108:29]
  wire [4:0] control_io_metadata_init_bits_desc_state_field_type_12_field_type; // @[FpgaCloudSerHw.scala 108:29]
  wire [15:0] control_io_metadata_init_bits_desc_state_field_type_12_sub_class_id; // @[FpgaCloudSerHw.scala 108:29]
  wire  control_io_metadata_init_bits_desc_state_field_type_12_is_host; // @[FpgaCloudSerHw.scala 108:29]
  wire  control_io_metadata_init_bits_desc_state_field_type_13_is_repeated; // @[FpgaCloudSerHw.scala 108:29]
  wire [4:0] control_io_metadata_init_bits_desc_state_field_type_13_field_type; // @[FpgaCloudSerHw.scala 108:29]
  wire [15:0] control_io_metadata_init_bits_desc_state_field_type_13_sub_class_id; // @[FpgaCloudSerHw.scala 108:29]
  wire  control_io_metadata_init_bits_desc_state_field_type_13_is_host; // @[FpgaCloudSerHw.scala 108:29]
  wire  control_io_metadata_init_bits_desc_state_field_type_14_is_repeated; // @[FpgaCloudSerHw.scala 108:29]
  wire [4:0] control_io_metadata_init_bits_desc_state_field_type_14_field_type; // @[FpgaCloudSerHw.scala 108:29]
  wire [15:0] control_io_metadata_init_bits_desc_state_field_type_14_sub_class_id; // @[FpgaCloudSerHw.scala 108:29]
  wire  control_io_metadata_init_bits_desc_state_field_type_14_is_host; // @[FpgaCloudSerHw.scala 108:29]
  wire  control_io_metadata_init_bits_desc_state_field_type_15_is_repeated; // @[FpgaCloudSerHw.scala 108:29]
  wire [4:0] control_io_metadata_init_bits_desc_state_field_type_15_field_type; // @[FpgaCloudSerHw.scala 108:29]
  wire [15:0] control_io_metadata_init_bits_desc_state_field_type_15_sub_class_id; // @[FpgaCloudSerHw.scala 108:29]
  wire  control_io_metadata_init_bits_desc_state_field_type_15_is_host; // @[FpgaCloudSerHw.scala 108:29]
  wire  control_io_metadata_init_bits_desc_state_field_type_16_is_repeated; // @[FpgaCloudSerHw.scala 108:29]
  wire [4:0] control_io_metadata_init_bits_desc_state_field_type_16_field_type; // @[FpgaCloudSerHw.scala 108:29]
  wire [15:0] control_io_metadata_init_bits_desc_state_field_type_16_sub_class_id; // @[FpgaCloudSerHw.scala 108:29]
  wire  control_io_metadata_init_bits_desc_state_field_type_16_is_host; // @[FpgaCloudSerHw.scala 108:29]
  wire  control_io_metadata_init_bits_desc_state_field_type_17_is_repeated; // @[FpgaCloudSerHw.scala 108:29]
  wire [4:0] control_io_metadata_init_bits_desc_state_field_type_17_field_type; // @[FpgaCloudSerHw.scala 108:29]
  wire [15:0] control_io_metadata_init_bits_desc_state_field_type_17_sub_class_id; // @[FpgaCloudSerHw.scala 108:29]
  wire  control_io_metadata_init_bits_desc_state_field_type_17_is_host; // @[FpgaCloudSerHw.scala 108:29]
  wire  control_io_metadata_init_bits_desc_state_field_type_18_is_repeated; // @[FpgaCloudSerHw.scala 108:29]
  wire [4:0] control_io_metadata_init_bits_desc_state_field_type_18_field_type; // @[FpgaCloudSerHw.scala 108:29]
  wire [15:0] control_io_metadata_init_bits_desc_state_field_type_18_sub_class_id; // @[FpgaCloudSerHw.scala 108:29]
  wire  control_io_metadata_init_bits_desc_state_field_type_18_is_host; // @[FpgaCloudSerHw.scala 108:29]
  wire  control_io_metadata_init_bits_desc_state_field_type_19_is_repeated; // @[FpgaCloudSerHw.scala 108:29]
  wire [4:0] control_io_metadata_init_bits_desc_state_field_type_19_field_type; // @[FpgaCloudSerHw.scala 108:29]
  wire [15:0] control_io_metadata_init_bits_desc_state_field_type_19_sub_class_id; // @[FpgaCloudSerHw.scala 108:29]
  wire  control_io_metadata_init_bits_desc_state_field_type_19_is_host; // @[FpgaCloudSerHw.scala 108:29]
  wire  control_io_metadata_init_bits_desc_state_field_type_20_is_repeated; // @[FpgaCloudSerHw.scala 108:29]
  wire [4:0] control_io_metadata_init_bits_desc_state_field_type_20_field_type; // @[FpgaCloudSerHw.scala 108:29]
  wire [15:0] control_io_metadata_init_bits_desc_state_field_type_20_sub_class_id; // @[FpgaCloudSerHw.scala 108:29]
  wire  control_io_metadata_init_bits_desc_state_field_type_20_is_host; // @[FpgaCloudSerHw.scala 108:29]
  wire  control_io_metadata_init_bits_desc_state_field_type_21_is_repeated; // @[FpgaCloudSerHw.scala 108:29]
  wire [4:0] control_io_metadata_init_bits_desc_state_field_type_21_field_type; // @[FpgaCloudSerHw.scala 108:29]
  wire [15:0] control_io_metadata_init_bits_desc_state_field_type_21_sub_class_id; // @[FpgaCloudSerHw.scala 108:29]
  wire  control_io_metadata_init_bits_desc_state_field_type_21_is_host; // @[FpgaCloudSerHw.scala 108:29]
  wire  control_io_metadata_init_bits_desc_state_field_type_22_is_repeated; // @[FpgaCloudSerHw.scala 108:29]
  wire [4:0] control_io_metadata_init_bits_desc_state_field_type_22_field_type; // @[FpgaCloudSerHw.scala 108:29]
  wire [15:0] control_io_metadata_init_bits_desc_state_field_type_22_sub_class_id; // @[FpgaCloudSerHw.scala 108:29]
  wire  control_io_metadata_init_bits_desc_state_field_type_22_is_host; // @[FpgaCloudSerHw.scala 108:29]
  wire  control_io_metadata_init_bits_desc_state_field_type_23_is_repeated; // @[FpgaCloudSerHw.scala 108:29]
  wire [4:0] control_io_metadata_init_bits_desc_state_field_type_23_field_type; // @[FpgaCloudSerHw.scala 108:29]
  wire [15:0] control_io_metadata_init_bits_desc_state_field_type_23_sub_class_id; // @[FpgaCloudSerHw.scala 108:29]
  wire  control_io_metadata_init_bits_desc_state_field_type_23_is_host; // @[FpgaCloudSerHw.scala 108:29]
  wire  control_io_metadata_init_bits_desc_state_field_type_24_is_repeated; // @[FpgaCloudSerHw.scala 108:29]
  wire [4:0] control_io_metadata_init_bits_desc_state_field_type_24_field_type; // @[FpgaCloudSerHw.scala 108:29]
  wire [15:0] control_io_metadata_init_bits_desc_state_field_type_24_sub_class_id; // @[FpgaCloudSerHw.scala 108:29]
  wire  control_io_metadata_init_bits_desc_state_field_type_24_is_host; // @[FpgaCloudSerHw.scala 108:29]
  wire  control_io_metadata_init_bits_desc_state_field_type_25_is_repeated; // @[FpgaCloudSerHw.scala 108:29]
  wire [4:0] control_io_metadata_init_bits_desc_state_field_type_25_field_type; // @[FpgaCloudSerHw.scala 108:29]
  wire [15:0] control_io_metadata_init_bits_desc_state_field_type_25_sub_class_id; // @[FpgaCloudSerHw.scala 108:29]
  wire  control_io_metadata_init_bits_desc_state_field_type_25_is_host; // @[FpgaCloudSerHw.scala 108:29]
  wire  control_io_metadata_init_bits_desc_state_field_type_26_is_repeated; // @[FpgaCloudSerHw.scala 108:29]
  wire [4:0] control_io_metadata_init_bits_desc_state_field_type_26_field_type; // @[FpgaCloudSerHw.scala 108:29]
  wire [15:0] control_io_metadata_init_bits_desc_state_field_type_26_sub_class_id; // @[FpgaCloudSerHw.scala 108:29]
  wire  control_io_metadata_init_bits_desc_state_field_type_26_is_host; // @[FpgaCloudSerHw.scala 108:29]
  wire  control_io_metadata_init_bits_desc_state_field_type_27_is_repeated; // @[FpgaCloudSerHw.scala 108:29]
  wire [4:0] control_io_metadata_init_bits_desc_state_field_type_27_field_type; // @[FpgaCloudSerHw.scala 108:29]
  wire [15:0] control_io_metadata_init_bits_desc_state_field_type_27_sub_class_id; // @[FpgaCloudSerHw.scala 108:29]
  wire  control_io_metadata_init_bits_desc_state_field_type_27_is_host; // @[FpgaCloudSerHw.scala 108:29]
  wire  control_io_metadata_init_bits_desc_state_field_type_28_is_repeated; // @[FpgaCloudSerHw.scala 108:29]
  wire [4:0] control_io_metadata_init_bits_desc_state_field_type_28_field_type; // @[FpgaCloudSerHw.scala 108:29]
  wire [15:0] control_io_metadata_init_bits_desc_state_field_type_28_sub_class_id; // @[FpgaCloudSerHw.scala 108:29]
  wire  control_io_metadata_init_bits_desc_state_field_type_28_is_host; // @[FpgaCloudSerHw.scala 108:29]
  wire  control_io_metadata_init_bits_desc_state_field_type_29_is_repeated; // @[FpgaCloudSerHw.scala 108:29]
  wire [4:0] control_io_metadata_init_bits_desc_state_field_type_29_field_type; // @[FpgaCloudSerHw.scala 108:29]
  wire [15:0] control_io_metadata_init_bits_desc_state_field_type_29_sub_class_id; // @[FpgaCloudSerHw.scala 108:29]
  wire  control_io_metadata_init_bits_desc_state_field_type_29_is_host; // @[FpgaCloudSerHw.scala 108:29]
  wire  control_io_metadata_init_bits_desc_state_field_type_30_is_repeated; // @[FpgaCloudSerHw.scala 108:29]
  wire [4:0] control_io_metadata_init_bits_desc_state_field_type_30_field_type; // @[FpgaCloudSerHw.scala 108:29]
  wire [15:0] control_io_metadata_init_bits_desc_state_field_type_30_sub_class_id; // @[FpgaCloudSerHw.scala 108:29]
  wire  control_io_metadata_init_bits_desc_state_field_type_30_is_host; // @[FpgaCloudSerHw.scala 108:29]
  wire  control_io_metadata_init_bits_desc_state_field_type_31_is_repeated; // @[FpgaCloudSerHw.scala 108:29]
  wire [4:0] control_io_metadata_init_bits_desc_state_field_type_31_field_type; // @[FpgaCloudSerHw.scala 108:29]
  wire [15:0] control_io_metadata_init_bits_desc_state_field_type_31_sub_class_id; // @[FpgaCloudSerHw.scala 108:29]
  wire  control_io_metadata_init_bits_desc_state_field_type_31_is_host; // @[FpgaCloudSerHw.scala 108:29]
  wire  control_io_metadata_init_bits_desc_state_field_type_32_is_repeated; // @[FpgaCloudSerHw.scala 108:29]
  wire [4:0] control_io_metadata_init_bits_desc_state_field_type_32_field_type; // @[FpgaCloudSerHw.scala 108:29]
  wire [15:0] control_io_metadata_init_bits_desc_state_field_type_32_sub_class_id; // @[FpgaCloudSerHw.scala 108:29]
  wire  control_io_metadata_init_bits_desc_state_field_type_32_is_host; // @[FpgaCloudSerHw.scala 108:29]
  wire  control_io_ser_cmd_ready; // @[FpgaCloudSerHw.scala 108:29]
  wire  control_io_ser_cmd_valid; // @[FpgaCloudSerHw.scala 108:29]
  wire [9:0] control_io_ser_cmd_bits_class_id; // @[FpgaCloudSerHw.scala 108:29]
  wire [63:0] control_io_ser_cmd_bits_host_base_addr; // @[FpgaCloudSerHw.scala 108:29]
  wire  instIlaDbg_clk; // @[FpgaCloudSerHw.scala 166:40]
  wire  instIlaDbg_data_1; // @[FpgaCloudSerHw.scala 166:40]
  wire [31:0] instIlaDbg_data_0; // @[FpgaCloudSerHw.scala 166:40]
  reg  hbmRstn; // @[FpgaCloudSerHw.scala 52:77]
  wire  userRstn = ~reset & ~qdma_io_reg_control_0[0]; // @[FpgaCloudSerHw.scala 83:74]
  wire  _T = ~userRstn; // @[FpgaCloudSerHw.scala 101:33]
  reg  timer_en; // @[FpgaCloudSerHw.scala 145:39]
  reg  done_en; // @[FpgaCloudSerHw.scala 146:38]
  reg [31:0] timer_cnt; // @[FpgaCloudSerHw.scala 147:40]
  wire  _T_1 = control_io_ser_cmd_ready & control_io_ser_cmd_valid; // @[Decoupled.scala 40:37]
  wire  _T_2 = ser_io_done_ready & ser_io_done_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_0 = _T_2 ? 1'h0 : timer_en; // @[FpgaCloudSerHw.scala 151:48 FpgaCloudSerHw.scala 152:41 FpgaCloudSerHw.scala 154:41]
  wire  _GEN_1 = _T_1 | _GEN_0; // @[FpgaCloudSerHw.scala 149:50 FpgaCloudSerHw.scala 150:41]
  wire [31:0] _timer_cnt_T_1 = timer_cnt + 32'h1; // @[FpgaCloudSerHw.scala 160:54]
  wire  _GEN_4 = _T_2 | done_en; // @[FpgaCloudSerHw.scala 174:48 FpgaCloudSerHw.scala 175:41 FpgaCloudSerHw.scala 177:33]
  wire  report_w1_1 = qdma_io_out_ready_0;
  wire  report_w1_0 = qdma_io_out_valid_1;
  wire  report_w1_3 = qdma_io_out_ready_1;
  wire  report_w1_2 = qdma_io_out_valid;
  wire  report_w1_5 = qdma_io_out_ready;
  wire  report_w1_4 = qdma_io_out_valid_0;
  wire  report_w1_7 = qdma_io_in_ready;
  wire  report_w1_6 = qdma_io_in_valid;
  wire [15:0] qdma_io_reg_status_414_lo = {8'h0,report_w1_7,report_w1_6,report_w1_5,report_w1_4,report_w1_3,report_w1_2,
    report_w1_1,report_w1_0}; // @[Collector.scala 237:73]
  DebugBridge dbgBridgeInst ( // @[DebugBridge.scala 58:37]
    .clk(dbgBridgeInst_clk),
    .S_BSCAN_drck(dbgBridgeInst_S_BSCAN_drck),
    .S_BSCAN_shift(dbgBridgeInst_S_BSCAN_shift),
    .S_BSCAN_tdi(dbgBridgeInst_S_BSCAN_tdi),
    .S_BSCAN_update(dbgBridgeInst_S_BSCAN_update),
    .S_BSCAN_sel(dbgBridgeInst_S_BSCAN_sel),
    .S_BSCAN_tdo(dbgBridgeInst_S_BSCAN_tdo),
    .S_BSCAN_tms(dbgBridgeInst_S_BSCAN_tms),
    .S_BSCAN_tck(dbgBridgeInst_S_BSCAN_tck),
    .S_BSCAN_runtest(dbgBridgeInst_S_BSCAN_runtest),
    .S_BSCAN_reset(dbgBridgeInst_S_BSCAN_reset),
    .S_BSCAN_capture(dbgBridgeInst_S_BSCAN_capture),
    .S_BSCAN_bscanid_en(dbgBridgeInst_S_BSCAN_bscanid_en)
  );
  HBM_DRIVER hbmDriver ( // @[FpgaCloudSerHw.scala 49:70]
    .clock(hbmDriver_clock),
    .io_hbm_clk(hbmDriver_io_hbm_clk),
    .io_hbm_rstn(hbmDriver_io_hbm_rstn)
  );
  QDMADynamic qdma ( // @[FpgaCloudSerHw.scala 68:26]
    .io_qdma_port_axi_aclk(qdma_io_qdma_port_axi_aclk),
    .io_qdma_port_axi_aresetn(qdma_io_qdma_port_axi_aresetn),
    .io_qdma_port_m_axib_awid(qdma_io_qdma_port_m_axib_awid),
    .io_qdma_port_m_axib_awaddr(qdma_io_qdma_port_m_axib_awaddr),
    .io_qdma_port_m_axib_awlen(qdma_io_qdma_port_m_axib_awlen),
    .io_qdma_port_m_axib_awsize(qdma_io_qdma_port_m_axib_awsize),
    .io_qdma_port_m_axib_awburst(qdma_io_qdma_port_m_axib_awburst),
    .io_qdma_port_m_axib_awprot(qdma_io_qdma_port_m_axib_awprot),
    .io_qdma_port_m_axib_awlock(qdma_io_qdma_port_m_axib_awlock),
    .io_qdma_port_m_axib_awcache(qdma_io_qdma_port_m_axib_awcache),
    .io_qdma_port_m_axib_awvalid(qdma_io_qdma_port_m_axib_awvalid),
    .io_qdma_port_m_axib_awready(qdma_io_qdma_port_m_axib_awready),
    .io_qdma_port_m_axib_wdata(qdma_io_qdma_port_m_axib_wdata),
    .io_qdma_port_m_axib_wstrb(qdma_io_qdma_port_m_axib_wstrb),
    .io_qdma_port_m_axib_wlast(qdma_io_qdma_port_m_axib_wlast),
    .io_qdma_port_m_axib_wvalid(qdma_io_qdma_port_m_axib_wvalid),
    .io_qdma_port_m_axib_wready(qdma_io_qdma_port_m_axib_wready),
    .io_qdma_port_m_axib_bid(qdma_io_qdma_port_m_axib_bid),
    .io_qdma_port_m_axib_bresp(qdma_io_qdma_port_m_axib_bresp),
    .io_qdma_port_m_axib_bvalid(qdma_io_qdma_port_m_axib_bvalid),
    .io_qdma_port_m_axib_bready(qdma_io_qdma_port_m_axib_bready),
    .io_qdma_port_m_axib_arid(qdma_io_qdma_port_m_axib_arid),
    .io_qdma_port_m_axib_araddr(qdma_io_qdma_port_m_axib_araddr),
    .io_qdma_port_m_axib_arlen(qdma_io_qdma_port_m_axib_arlen),
    .io_qdma_port_m_axib_arsize(qdma_io_qdma_port_m_axib_arsize),
    .io_qdma_port_m_axib_arburst(qdma_io_qdma_port_m_axib_arburst),
    .io_qdma_port_m_axib_arprot(qdma_io_qdma_port_m_axib_arprot),
    .io_qdma_port_m_axib_arlock(qdma_io_qdma_port_m_axib_arlock),
    .io_qdma_port_m_axib_arcache(qdma_io_qdma_port_m_axib_arcache),
    .io_qdma_port_m_axib_arvalid(qdma_io_qdma_port_m_axib_arvalid),
    .io_qdma_port_m_axib_arready(qdma_io_qdma_port_m_axib_arready),
    .io_qdma_port_m_axib_rid(qdma_io_qdma_port_m_axib_rid),
    .io_qdma_port_m_axib_rdata(qdma_io_qdma_port_m_axib_rdata),
    .io_qdma_port_m_axib_rresp(qdma_io_qdma_port_m_axib_rresp),
    .io_qdma_port_m_axib_rlast(qdma_io_qdma_port_m_axib_rlast),
    .io_qdma_port_m_axib_rvalid(qdma_io_qdma_port_m_axib_rvalid),
    .io_qdma_port_m_axib_rready(qdma_io_qdma_port_m_axib_rready),
    .io_qdma_port_m_axil_awaddr(qdma_io_qdma_port_m_axil_awaddr),
    .io_qdma_port_m_axil_awvalid(qdma_io_qdma_port_m_axil_awvalid),
    .io_qdma_port_m_axil_awready(qdma_io_qdma_port_m_axil_awready),
    .io_qdma_port_m_axil_wdata(qdma_io_qdma_port_m_axil_wdata),
    .io_qdma_port_m_axil_wstrb(qdma_io_qdma_port_m_axil_wstrb),
    .io_qdma_port_m_axil_wvalid(qdma_io_qdma_port_m_axil_wvalid),
    .io_qdma_port_m_axil_wready(qdma_io_qdma_port_m_axil_wready),
    .io_qdma_port_m_axil_bresp(qdma_io_qdma_port_m_axil_bresp),
    .io_qdma_port_m_axil_bvalid(qdma_io_qdma_port_m_axil_bvalid),
    .io_qdma_port_m_axil_bready(qdma_io_qdma_port_m_axil_bready),
    .io_qdma_port_m_axil_araddr(qdma_io_qdma_port_m_axil_araddr),
    .io_qdma_port_m_axil_arvalid(qdma_io_qdma_port_m_axil_arvalid),
    .io_qdma_port_m_axil_arready(qdma_io_qdma_port_m_axil_arready),
    .io_qdma_port_m_axil_rdata(qdma_io_qdma_port_m_axil_rdata),
    .io_qdma_port_m_axil_rresp(qdma_io_qdma_port_m_axil_rresp),
    .io_qdma_port_m_axil_rvalid(qdma_io_qdma_port_m_axil_rvalid),
    .io_qdma_port_m_axil_rready(qdma_io_qdma_port_m_axil_rready),
    .io_qdma_port_h2c_byp_in_st_addr(qdma_io_qdma_port_h2c_byp_in_st_addr),
    .io_qdma_port_h2c_byp_in_st_len(qdma_io_qdma_port_h2c_byp_in_st_len),
    .io_qdma_port_h2c_byp_in_st_eop(qdma_io_qdma_port_h2c_byp_in_st_eop),
    .io_qdma_port_h2c_byp_in_st_sop(qdma_io_qdma_port_h2c_byp_in_st_sop),
    .io_qdma_port_h2c_byp_in_st_mrkr_req(qdma_io_qdma_port_h2c_byp_in_st_mrkr_req),
    .io_qdma_port_h2c_byp_in_st_sdi(qdma_io_qdma_port_h2c_byp_in_st_sdi),
    .io_qdma_port_h2c_byp_in_st_qid(qdma_io_qdma_port_h2c_byp_in_st_qid),
    .io_qdma_port_h2c_byp_in_st_error(qdma_io_qdma_port_h2c_byp_in_st_error),
    .io_qdma_port_h2c_byp_in_st_func(qdma_io_qdma_port_h2c_byp_in_st_func),
    .io_qdma_port_h2c_byp_in_st_cidx(qdma_io_qdma_port_h2c_byp_in_st_cidx),
    .io_qdma_port_h2c_byp_in_st_port_id(qdma_io_qdma_port_h2c_byp_in_st_port_id),
    .io_qdma_port_h2c_byp_in_st_no_dma(qdma_io_qdma_port_h2c_byp_in_st_no_dma),
    .io_qdma_port_h2c_byp_in_st_vld(qdma_io_qdma_port_h2c_byp_in_st_vld),
    .io_qdma_port_h2c_byp_in_st_rdy(qdma_io_qdma_port_h2c_byp_in_st_rdy),
    .io_qdma_port_c2h_byp_in_st_csh_addr(qdma_io_qdma_port_c2h_byp_in_st_csh_addr),
    .io_qdma_port_c2h_byp_in_st_csh_qid(qdma_io_qdma_port_c2h_byp_in_st_csh_qid),
    .io_qdma_port_c2h_byp_in_st_csh_error(qdma_io_qdma_port_c2h_byp_in_st_csh_error),
    .io_qdma_port_c2h_byp_in_st_csh_func(qdma_io_qdma_port_c2h_byp_in_st_csh_func),
    .io_qdma_port_c2h_byp_in_st_csh_port_id(qdma_io_qdma_port_c2h_byp_in_st_csh_port_id),
    .io_qdma_port_c2h_byp_in_st_csh_pfch_tag(qdma_io_qdma_port_c2h_byp_in_st_csh_pfch_tag),
    .io_qdma_port_c2h_byp_in_st_csh_vld(qdma_io_qdma_port_c2h_byp_in_st_csh_vld),
    .io_qdma_port_c2h_byp_in_st_csh_rdy(qdma_io_qdma_port_c2h_byp_in_st_csh_rdy),
    .io_qdma_port_s_axis_c2h_tdata(qdma_io_qdma_port_s_axis_c2h_tdata),
    .io_qdma_port_s_axis_c2h_tcrc(qdma_io_qdma_port_s_axis_c2h_tcrc),
    .io_qdma_port_s_axis_c2h_ctrl_marker(qdma_io_qdma_port_s_axis_c2h_ctrl_marker),
    .io_qdma_port_s_axis_c2h_ctrl_ecc(qdma_io_qdma_port_s_axis_c2h_ctrl_ecc),
    .io_qdma_port_s_axis_c2h_ctrl_len(qdma_io_qdma_port_s_axis_c2h_ctrl_len),
    .io_qdma_port_s_axis_c2h_ctrl_port_id(qdma_io_qdma_port_s_axis_c2h_ctrl_port_id),
    .io_qdma_port_s_axis_c2h_ctrl_qid(qdma_io_qdma_port_s_axis_c2h_ctrl_qid),
    .io_qdma_port_s_axis_c2h_ctrl_has_cmpt(qdma_io_qdma_port_s_axis_c2h_ctrl_has_cmpt),
    .io_qdma_port_s_axis_c2h_mty(qdma_io_qdma_port_s_axis_c2h_mty),
    .io_qdma_port_s_axis_c2h_tlast(qdma_io_qdma_port_s_axis_c2h_tlast),
    .io_qdma_port_s_axis_c2h_tvalid(qdma_io_qdma_port_s_axis_c2h_tvalid),
    .io_qdma_port_s_axis_c2h_tready(qdma_io_qdma_port_s_axis_c2h_tready),
    .io_qdma_port_m_axis_h2c_tdata(qdma_io_qdma_port_m_axis_h2c_tdata),
    .io_qdma_port_m_axis_h2c_tcrc(qdma_io_qdma_port_m_axis_h2c_tcrc),
    .io_qdma_port_m_axis_h2c_tuser_qid(qdma_io_qdma_port_m_axis_h2c_tuser_qid),
    .io_qdma_port_m_axis_h2c_tuser_port_id(qdma_io_qdma_port_m_axis_h2c_tuser_port_id),
    .io_qdma_port_m_axis_h2c_tuser_err(qdma_io_qdma_port_m_axis_h2c_tuser_err),
    .io_qdma_port_m_axis_h2c_tuser_mdata(qdma_io_qdma_port_m_axis_h2c_tuser_mdata),
    .io_qdma_port_m_axis_h2c_tuser_mty(qdma_io_qdma_port_m_axis_h2c_tuser_mty),
    .io_qdma_port_m_axis_h2c_tuser_zero_byte(qdma_io_qdma_port_m_axis_h2c_tuser_zero_byte),
    .io_qdma_port_m_axis_h2c_tlast(qdma_io_qdma_port_m_axis_h2c_tlast),
    .io_qdma_port_m_axis_h2c_tvalid(qdma_io_qdma_port_m_axis_h2c_tvalid),
    .io_qdma_port_m_axis_h2c_tready(qdma_io_qdma_port_m_axis_h2c_tready),
    .io_user_clk(qdma_io_user_clk),
    .io_user_arstn(qdma_io_user_arstn),
    .io_h2c_cmd_ready(qdma_io_h2c_cmd_ready),
    .io_h2c_cmd_valid(qdma_io_h2c_cmd_valid),
    .io_h2c_cmd_bits_addr(qdma_io_h2c_cmd_bits_addr),
    .io_h2c_cmd_bits_len(qdma_io_h2c_cmd_bits_len),
    .io_h2c_data_valid(qdma_io_h2c_data_valid),
    .io_reg_control_0(qdma_io_reg_control_0),
    .io_reg_control_8(qdma_io_reg_control_8),
    .io_reg_control_9(qdma_io_reg_control_9),
    .io_reg_control_10(qdma_io_reg_control_10),
    .io_reg_control_11(qdma_io_reg_control_11),
    .io_reg_control_12(qdma_io_reg_control_12),
    .io_reg_control_13(qdma_io_reg_control_13),
    .io_reg_control_14(qdma_io_reg_control_14),
    .io_reg_status_300(qdma_io_reg_status_300),
    .io_reg_status_400(qdma_io_reg_status_400),
    .io_reg_status_401(qdma_io_reg_status_401),
    .io_reg_status_402(qdma_io_reg_status_402),
    .io_reg_status_403(qdma_io_reg_status_403),
    .io_reg_status_404(qdma_io_reg_status_404),
    .io_reg_status_405(qdma_io_reg_status_405),
    .io_reg_status_406(qdma_io_reg_status_406),
    .io_reg_status_407(qdma_io_reg_status_407),
    .io_reg_status_408(qdma_io_reg_status_408),
    .io_reg_status_409(qdma_io_reg_status_409),
    .io_reg_status_410(qdma_io_reg_status_410),
    .io_reg_status_411(qdma_io_reg_status_411),
    .io_reg_status_412(qdma_io_reg_status_412),
    .io_reg_status_413(qdma_io_reg_status_413),
    .io_reg_status_414(qdma_io_reg_status_414),
    .io_axib_aw_ready(qdma_io_axib_aw_ready),
    .io_axib_aw_valid(qdma_io_axib_aw_valid),
    .io_axib_aw_bits_addr(qdma_io_axib_aw_bits_addr),
    .io_axib_w_ready(qdma_io_axib_w_ready),
    .io_axib_w_valid(qdma_io_axib_w_valid),
    .io_axib_w_bits_data(qdma_io_axib_w_bits_data),
    .io_axib_r_ready(qdma_io_axib_r_ready),
    .io_axib_r_bits_data(qdma_io_axib_r_bits_data),
    .io_out_valid(qdma_io_out_valid),
    .counter_4_0(qdma_counter_4_0),
    .io_out_ready(qdma_io_out_ready),
    .counter_7_0(qdma_counter_7_0),
    .counter_1_0(qdma_counter_1_0),
    .io_in_ready(qdma_io_in_ready),
    .counter_3_1(qdma_counter_3_1),
    .io_out_ready_0(qdma_io_out_ready_0),
    .counter_6_0(qdma_counter_6_0),
    .io_out_valid_0(qdma_io_out_valid_0),
    .counter_0(qdma_counter_0),
    .io_in_valid(qdma_io_in_valid),
    .io_tlb_miss_count(qdma_io_tlb_miss_count),
    .io_out_valid_1(qdma_io_out_valid_1),
    .counter_2_1(qdma_counter_2_1),
    .counter_5_0(qdma_counter_5_0),
    .io_out_ready_1(qdma_io_out_ready_1)
  );
  Serializerhw ser ( // @[FpgaCloudSerHw.scala 104:21]
    .clock(ser_clock),
    .reset(ser_reset),
    .io_meta_in_ready(ser_io_meta_in_ready),
    .io_meta_in_valid(ser_io_meta_in_valid),
    .io_meta_in_bits_class_id(ser_io_meta_in_bits_class_id),
    .io_meta_in_bits_host_base_addr(ser_io_meta_in_bits_host_base_addr),
    .io_host_data_in_ready(ser_io_host_data_in_ready),
    .io_host_data_in_valid(ser_io_host_data_in_valid),
    .io_host_data_cmd_ready(ser_io_host_data_cmd_ready),
    .io_host_data_cmd_valid(ser_io_host_data_cmd_valid),
    .io_host_data_cmd_bits_vaddr(ser_io_host_data_cmd_bits_vaddr),
    .io_host_data_cmd_bits_length(ser_io_host_data_cmd_bits_length),
    .io_class_meta_req_ready(ser_io_class_meta_req_ready),
    .io_class_meta_req_valid(ser_io_class_meta_req_valid),
    .io_class_meta_req_bits_class_id(ser_io_class_meta_req_bits_class_id),
    .io_class_meta_rsp_valid(ser_io_class_meta_rsp_valid),
    .io_class_meta_rsp_bits_class_meta_max_field_num(ser_io_class_meta_rsp_bits_class_meta_max_field_num),
    .io_class_meta_rsp_bits_class_meta_field_type_0_is_repeated(
      ser_io_class_meta_rsp_bits_class_meta_field_type_0_is_repeated),
    .io_class_meta_rsp_bits_class_meta_field_type_0_field_type(
      ser_io_class_meta_rsp_bits_class_meta_field_type_0_field_type),
    .io_class_meta_rsp_bits_class_meta_field_type_0_sub_class_id(
      ser_io_class_meta_rsp_bits_class_meta_field_type_0_sub_class_id),
    .io_class_meta_rsp_bits_class_meta_field_type_1_is_repeated(
      ser_io_class_meta_rsp_bits_class_meta_field_type_1_is_repeated),
    .io_class_meta_rsp_bits_class_meta_field_type_1_field_type(
      ser_io_class_meta_rsp_bits_class_meta_field_type_1_field_type),
    .io_class_meta_rsp_bits_class_meta_field_type_1_sub_class_id(
      ser_io_class_meta_rsp_bits_class_meta_field_type_1_sub_class_id),
    .io_class_meta_rsp_bits_class_meta_field_type_2_is_repeated(
      ser_io_class_meta_rsp_bits_class_meta_field_type_2_is_repeated),
    .io_class_meta_rsp_bits_class_meta_field_type_2_field_type(
      ser_io_class_meta_rsp_bits_class_meta_field_type_2_field_type),
    .io_class_meta_rsp_bits_class_meta_field_type_2_sub_class_id(
      ser_io_class_meta_rsp_bits_class_meta_field_type_2_sub_class_id),
    .io_class_meta_rsp_bits_class_meta_field_type_3_is_repeated(
      ser_io_class_meta_rsp_bits_class_meta_field_type_3_is_repeated),
    .io_class_meta_rsp_bits_class_meta_field_type_3_field_type(
      ser_io_class_meta_rsp_bits_class_meta_field_type_3_field_type),
    .io_class_meta_rsp_bits_class_meta_field_type_3_sub_class_id(
      ser_io_class_meta_rsp_bits_class_meta_field_type_3_sub_class_id),
    .io_class_meta_rsp_bits_class_meta_field_type_4_is_repeated(
      ser_io_class_meta_rsp_bits_class_meta_field_type_4_is_repeated),
    .io_class_meta_rsp_bits_class_meta_field_type_4_field_type(
      ser_io_class_meta_rsp_bits_class_meta_field_type_4_field_type),
    .io_class_meta_rsp_bits_class_meta_field_type_4_sub_class_id(
      ser_io_class_meta_rsp_bits_class_meta_field_type_4_sub_class_id),
    .io_class_meta_rsp_bits_class_meta_field_type_5_is_repeated(
      ser_io_class_meta_rsp_bits_class_meta_field_type_5_is_repeated),
    .io_class_meta_rsp_bits_class_meta_field_type_5_field_type(
      ser_io_class_meta_rsp_bits_class_meta_field_type_5_field_type),
    .io_class_meta_rsp_bits_class_meta_field_type_5_sub_class_id(
      ser_io_class_meta_rsp_bits_class_meta_field_type_5_sub_class_id),
    .io_class_meta_rsp_bits_class_meta_field_type_6_is_repeated(
      ser_io_class_meta_rsp_bits_class_meta_field_type_6_is_repeated),
    .io_class_meta_rsp_bits_class_meta_field_type_6_field_type(
      ser_io_class_meta_rsp_bits_class_meta_field_type_6_field_type),
    .io_class_meta_rsp_bits_class_meta_field_type_6_sub_class_id(
      ser_io_class_meta_rsp_bits_class_meta_field_type_6_sub_class_id),
    .io_class_meta_rsp_bits_class_meta_field_type_7_is_repeated(
      ser_io_class_meta_rsp_bits_class_meta_field_type_7_is_repeated),
    .io_class_meta_rsp_bits_class_meta_field_type_7_field_type(
      ser_io_class_meta_rsp_bits_class_meta_field_type_7_field_type),
    .io_class_meta_rsp_bits_class_meta_field_type_7_sub_class_id(
      ser_io_class_meta_rsp_bits_class_meta_field_type_7_sub_class_id),
    .io_class_meta_rsp_bits_class_meta_field_type_8_is_repeated(
      ser_io_class_meta_rsp_bits_class_meta_field_type_8_is_repeated),
    .io_class_meta_rsp_bits_class_meta_field_type_8_field_type(
      ser_io_class_meta_rsp_bits_class_meta_field_type_8_field_type),
    .io_class_meta_rsp_bits_class_meta_field_type_8_sub_class_id(
      ser_io_class_meta_rsp_bits_class_meta_field_type_8_sub_class_id),
    .io_class_meta_rsp_bits_class_meta_field_type_9_is_repeated(
      ser_io_class_meta_rsp_bits_class_meta_field_type_9_is_repeated),
    .io_class_meta_rsp_bits_class_meta_field_type_9_field_type(
      ser_io_class_meta_rsp_bits_class_meta_field_type_9_field_type),
    .io_class_meta_rsp_bits_class_meta_field_type_9_sub_class_id(
      ser_io_class_meta_rsp_bits_class_meta_field_type_9_sub_class_id),
    .io_class_meta_rsp_bits_class_meta_field_type_10_is_repeated(
      ser_io_class_meta_rsp_bits_class_meta_field_type_10_is_repeated),
    .io_class_meta_rsp_bits_class_meta_field_type_10_field_type(
      ser_io_class_meta_rsp_bits_class_meta_field_type_10_field_type),
    .io_class_meta_rsp_bits_class_meta_field_type_10_sub_class_id(
      ser_io_class_meta_rsp_bits_class_meta_field_type_10_sub_class_id),
    .io_class_meta_rsp_bits_class_meta_field_type_11_is_repeated(
      ser_io_class_meta_rsp_bits_class_meta_field_type_11_is_repeated),
    .io_class_meta_rsp_bits_class_meta_field_type_11_field_type(
      ser_io_class_meta_rsp_bits_class_meta_field_type_11_field_type),
    .io_class_meta_rsp_bits_class_meta_field_type_11_sub_class_id(
      ser_io_class_meta_rsp_bits_class_meta_field_type_11_sub_class_id),
    .io_class_meta_rsp_bits_class_meta_field_type_12_is_repeated(
      ser_io_class_meta_rsp_bits_class_meta_field_type_12_is_repeated),
    .io_class_meta_rsp_bits_class_meta_field_type_12_field_type(
      ser_io_class_meta_rsp_bits_class_meta_field_type_12_field_type),
    .io_class_meta_rsp_bits_class_meta_field_type_12_sub_class_id(
      ser_io_class_meta_rsp_bits_class_meta_field_type_12_sub_class_id),
    .io_class_meta_rsp_bits_class_meta_field_type_13_is_repeated(
      ser_io_class_meta_rsp_bits_class_meta_field_type_13_is_repeated),
    .io_class_meta_rsp_bits_class_meta_field_type_13_field_type(
      ser_io_class_meta_rsp_bits_class_meta_field_type_13_field_type),
    .io_class_meta_rsp_bits_class_meta_field_type_13_sub_class_id(
      ser_io_class_meta_rsp_bits_class_meta_field_type_13_sub_class_id),
    .io_class_meta_rsp_bits_class_meta_field_type_14_is_repeated(
      ser_io_class_meta_rsp_bits_class_meta_field_type_14_is_repeated),
    .io_class_meta_rsp_bits_class_meta_field_type_14_field_type(
      ser_io_class_meta_rsp_bits_class_meta_field_type_14_field_type),
    .io_class_meta_rsp_bits_class_meta_field_type_14_sub_class_id(
      ser_io_class_meta_rsp_bits_class_meta_field_type_14_sub_class_id),
    .io_class_meta_rsp_bits_class_meta_field_type_15_is_repeated(
      ser_io_class_meta_rsp_bits_class_meta_field_type_15_is_repeated),
    .io_class_meta_rsp_bits_class_meta_field_type_15_field_type(
      ser_io_class_meta_rsp_bits_class_meta_field_type_15_field_type),
    .io_class_meta_rsp_bits_class_meta_field_type_15_sub_class_id(
      ser_io_class_meta_rsp_bits_class_meta_field_type_15_sub_class_id),
    .io_class_meta_rsp_bits_class_meta_field_type_16_is_repeated(
      ser_io_class_meta_rsp_bits_class_meta_field_type_16_is_repeated),
    .io_class_meta_rsp_bits_class_meta_field_type_16_field_type(
      ser_io_class_meta_rsp_bits_class_meta_field_type_16_field_type),
    .io_class_meta_rsp_bits_class_meta_field_type_16_sub_class_id(
      ser_io_class_meta_rsp_bits_class_meta_field_type_16_sub_class_id),
    .io_class_meta_rsp_bits_class_meta_field_type_17_is_repeated(
      ser_io_class_meta_rsp_bits_class_meta_field_type_17_is_repeated),
    .io_class_meta_rsp_bits_class_meta_field_type_17_field_type(
      ser_io_class_meta_rsp_bits_class_meta_field_type_17_field_type),
    .io_class_meta_rsp_bits_class_meta_field_type_17_sub_class_id(
      ser_io_class_meta_rsp_bits_class_meta_field_type_17_sub_class_id),
    .io_class_meta_rsp_bits_class_meta_field_type_18_is_repeated(
      ser_io_class_meta_rsp_bits_class_meta_field_type_18_is_repeated),
    .io_class_meta_rsp_bits_class_meta_field_type_18_field_type(
      ser_io_class_meta_rsp_bits_class_meta_field_type_18_field_type),
    .io_class_meta_rsp_bits_class_meta_field_type_18_sub_class_id(
      ser_io_class_meta_rsp_bits_class_meta_field_type_18_sub_class_id),
    .io_class_meta_rsp_bits_class_meta_field_type_19_is_repeated(
      ser_io_class_meta_rsp_bits_class_meta_field_type_19_is_repeated),
    .io_class_meta_rsp_bits_class_meta_field_type_19_field_type(
      ser_io_class_meta_rsp_bits_class_meta_field_type_19_field_type),
    .io_class_meta_rsp_bits_class_meta_field_type_19_sub_class_id(
      ser_io_class_meta_rsp_bits_class_meta_field_type_19_sub_class_id),
    .io_class_meta_rsp_bits_class_meta_field_type_20_is_repeated(
      ser_io_class_meta_rsp_bits_class_meta_field_type_20_is_repeated),
    .io_class_meta_rsp_bits_class_meta_field_type_20_field_type(
      ser_io_class_meta_rsp_bits_class_meta_field_type_20_field_type),
    .io_class_meta_rsp_bits_class_meta_field_type_20_sub_class_id(
      ser_io_class_meta_rsp_bits_class_meta_field_type_20_sub_class_id),
    .io_class_meta_rsp_bits_class_meta_field_type_21_is_repeated(
      ser_io_class_meta_rsp_bits_class_meta_field_type_21_is_repeated),
    .io_class_meta_rsp_bits_class_meta_field_type_21_field_type(
      ser_io_class_meta_rsp_bits_class_meta_field_type_21_field_type),
    .io_class_meta_rsp_bits_class_meta_field_type_21_sub_class_id(
      ser_io_class_meta_rsp_bits_class_meta_field_type_21_sub_class_id),
    .io_class_meta_rsp_bits_class_meta_field_type_22_is_repeated(
      ser_io_class_meta_rsp_bits_class_meta_field_type_22_is_repeated),
    .io_class_meta_rsp_bits_class_meta_field_type_22_field_type(
      ser_io_class_meta_rsp_bits_class_meta_field_type_22_field_type),
    .io_class_meta_rsp_bits_class_meta_field_type_22_sub_class_id(
      ser_io_class_meta_rsp_bits_class_meta_field_type_22_sub_class_id),
    .io_class_meta_rsp_bits_class_meta_field_type_23_is_repeated(
      ser_io_class_meta_rsp_bits_class_meta_field_type_23_is_repeated),
    .io_class_meta_rsp_bits_class_meta_field_type_23_field_type(
      ser_io_class_meta_rsp_bits_class_meta_field_type_23_field_type),
    .io_class_meta_rsp_bits_class_meta_field_type_23_sub_class_id(
      ser_io_class_meta_rsp_bits_class_meta_field_type_23_sub_class_id),
    .io_class_meta_rsp_bits_class_meta_field_type_24_is_repeated(
      ser_io_class_meta_rsp_bits_class_meta_field_type_24_is_repeated),
    .io_class_meta_rsp_bits_class_meta_field_type_24_field_type(
      ser_io_class_meta_rsp_bits_class_meta_field_type_24_field_type),
    .io_class_meta_rsp_bits_class_meta_field_type_24_sub_class_id(
      ser_io_class_meta_rsp_bits_class_meta_field_type_24_sub_class_id),
    .io_class_meta_rsp_bits_class_meta_field_type_25_is_repeated(
      ser_io_class_meta_rsp_bits_class_meta_field_type_25_is_repeated),
    .io_class_meta_rsp_bits_class_meta_field_type_25_field_type(
      ser_io_class_meta_rsp_bits_class_meta_field_type_25_field_type),
    .io_class_meta_rsp_bits_class_meta_field_type_25_sub_class_id(
      ser_io_class_meta_rsp_bits_class_meta_field_type_25_sub_class_id),
    .io_class_meta_rsp_bits_class_meta_field_type_26_is_repeated(
      ser_io_class_meta_rsp_bits_class_meta_field_type_26_is_repeated),
    .io_class_meta_rsp_bits_class_meta_field_type_26_field_type(
      ser_io_class_meta_rsp_bits_class_meta_field_type_26_field_type),
    .io_class_meta_rsp_bits_class_meta_field_type_26_sub_class_id(
      ser_io_class_meta_rsp_bits_class_meta_field_type_26_sub_class_id),
    .io_class_meta_rsp_bits_class_meta_field_type_27_is_repeated(
      ser_io_class_meta_rsp_bits_class_meta_field_type_27_is_repeated),
    .io_class_meta_rsp_bits_class_meta_field_type_27_field_type(
      ser_io_class_meta_rsp_bits_class_meta_field_type_27_field_type),
    .io_class_meta_rsp_bits_class_meta_field_type_27_sub_class_id(
      ser_io_class_meta_rsp_bits_class_meta_field_type_27_sub_class_id),
    .io_class_meta_rsp_bits_class_meta_field_type_28_is_repeated(
      ser_io_class_meta_rsp_bits_class_meta_field_type_28_is_repeated),
    .io_class_meta_rsp_bits_class_meta_field_type_28_field_type(
      ser_io_class_meta_rsp_bits_class_meta_field_type_28_field_type),
    .io_class_meta_rsp_bits_class_meta_field_type_28_sub_class_id(
      ser_io_class_meta_rsp_bits_class_meta_field_type_28_sub_class_id),
    .io_class_meta_rsp_bits_class_meta_field_type_29_is_repeated(
      ser_io_class_meta_rsp_bits_class_meta_field_type_29_is_repeated),
    .io_class_meta_rsp_bits_class_meta_field_type_29_field_type(
      ser_io_class_meta_rsp_bits_class_meta_field_type_29_field_type),
    .io_class_meta_rsp_bits_class_meta_field_type_29_sub_class_id(
      ser_io_class_meta_rsp_bits_class_meta_field_type_29_sub_class_id),
    .io_class_meta_rsp_bits_class_meta_field_type_30_is_repeated(
      ser_io_class_meta_rsp_bits_class_meta_field_type_30_is_repeated),
    .io_class_meta_rsp_bits_class_meta_field_type_30_field_type(
      ser_io_class_meta_rsp_bits_class_meta_field_type_30_field_type),
    .io_class_meta_rsp_bits_class_meta_field_type_30_sub_class_id(
      ser_io_class_meta_rsp_bits_class_meta_field_type_30_sub_class_id),
    .io_class_meta_rsp_bits_class_meta_field_type_31_is_repeated(
      ser_io_class_meta_rsp_bits_class_meta_field_type_31_is_repeated),
    .io_class_meta_rsp_bits_class_meta_field_type_31_field_type(
      ser_io_class_meta_rsp_bits_class_meta_field_type_31_field_type),
    .io_class_meta_rsp_bits_class_meta_field_type_31_sub_class_id(
      ser_io_class_meta_rsp_bits_class_meta_field_type_31_sub_class_id),
    .io_class_meta_rsp_bits_class_meta_field_type_32_is_repeated(
      ser_io_class_meta_rsp_bits_class_meta_field_type_32_is_repeated),
    .io_class_meta_rsp_bits_class_meta_field_type_32_field_type(
      ser_io_class_meta_rsp_bits_class_meta_field_type_32_field_type),
    .io_class_meta_rsp_bits_class_meta_field_type_32_sub_class_id(
      ser_io_class_meta_rsp_bits_class_meta_field_type_32_sub_class_id),
    .io_done_ready(ser_io_done_ready),
    .io_done_valid(ser_io_done_valid),
    .counter_3_0(ser_counter_3_0),
    .counter_2_0(ser_counter_2_0),
    .counter_8(ser_counter_8),
    .counter_1_1(ser_counter_1_1)
  );
  ClassMetaTable meta_table ( // @[FpgaCloudSerHw.scala 105:28]
    .clock(meta_table_clock),
    .reset(meta_table_reset),
    .io_class_meta_init_ready(meta_table_io_class_meta_init_ready),
    .io_class_meta_init_valid(meta_table_io_class_meta_init_valid),
    .io_class_meta_init_bits_class_id(meta_table_io_class_meta_init_bits_class_id),
    .io_class_meta_init_bits_desc_state_class_length(meta_table_io_class_meta_init_bits_desc_state_class_length),
    .io_class_meta_init_bits_desc_state_max_field_num(meta_table_io_class_meta_init_bits_desc_state_max_field_num),
    .io_class_meta_init_bits_desc_state_field_type_0_is_repeated(
      meta_table_io_class_meta_init_bits_desc_state_field_type_0_is_repeated),
    .io_class_meta_init_bits_desc_state_field_type_0_field_type(
      meta_table_io_class_meta_init_bits_desc_state_field_type_0_field_type),
    .io_class_meta_init_bits_desc_state_field_type_0_sub_class_id(
      meta_table_io_class_meta_init_bits_desc_state_field_type_0_sub_class_id),
    .io_class_meta_init_bits_desc_state_field_type_0_is_host(
      meta_table_io_class_meta_init_bits_desc_state_field_type_0_is_host),
    .io_class_meta_init_bits_desc_state_field_type_1_is_repeated(
      meta_table_io_class_meta_init_bits_desc_state_field_type_1_is_repeated),
    .io_class_meta_init_bits_desc_state_field_type_1_field_type(
      meta_table_io_class_meta_init_bits_desc_state_field_type_1_field_type),
    .io_class_meta_init_bits_desc_state_field_type_1_sub_class_id(
      meta_table_io_class_meta_init_bits_desc_state_field_type_1_sub_class_id),
    .io_class_meta_init_bits_desc_state_field_type_1_is_host(
      meta_table_io_class_meta_init_bits_desc_state_field_type_1_is_host),
    .io_class_meta_init_bits_desc_state_field_type_2_is_repeated(
      meta_table_io_class_meta_init_bits_desc_state_field_type_2_is_repeated),
    .io_class_meta_init_bits_desc_state_field_type_2_field_type(
      meta_table_io_class_meta_init_bits_desc_state_field_type_2_field_type),
    .io_class_meta_init_bits_desc_state_field_type_2_sub_class_id(
      meta_table_io_class_meta_init_bits_desc_state_field_type_2_sub_class_id),
    .io_class_meta_init_bits_desc_state_field_type_2_is_host(
      meta_table_io_class_meta_init_bits_desc_state_field_type_2_is_host),
    .io_class_meta_init_bits_desc_state_field_type_3_is_repeated(
      meta_table_io_class_meta_init_bits_desc_state_field_type_3_is_repeated),
    .io_class_meta_init_bits_desc_state_field_type_3_field_type(
      meta_table_io_class_meta_init_bits_desc_state_field_type_3_field_type),
    .io_class_meta_init_bits_desc_state_field_type_3_sub_class_id(
      meta_table_io_class_meta_init_bits_desc_state_field_type_3_sub_class_id),
    .io_class_meta_init_bits_desc_state_field_type_3_is_host(
      meta_table_io_class_meta_init_bits_desc_state_field_type_3_is_host),
    .io_class_meta_init_bits_desc_state_field_type_4_is_repeated(
      meta_table_io_class_meta_init_bits_desc_state_field_type_4_is_repeated),
    .io_class_meta_init_bits_desc_state_field_type_4_field_type(
      meta_table_io_class_meta_init_bits_desc_state_field_type_4_field_type),
    .io_class_meta_init_bits_desc_state_field_type_4_sub_class_id(
      meta_table_io_class_meta_init_bits_desc_state_field_type_4_sub_class_id),
    .io_class_meta_init_bits_desc_state_field_type_4_is_host(
      meta_table_io_class_meta_init_bits_desc_state_field_type_4_is_host),
    .io_class_meta_init_bits_desc_state_field_type_5_is_repeated(
      meta_table_io_class_meta_init_bits_desc_state_field_type_5_is_repeated),
    .io_class_meta_init_bits_desc_state_field_type_5_field_type(
      meta_table_io_class_meta_init_bits_desc_state_field_type_5_field_type),
    .io_class_meta_init_bits_desc_state_field_type_5_sub_class_id(
      meta_table_io_class_meta_init_bits_desc_state_field_type_5_sub_class_id),
    .io_class_meta_init_bits_desc_state_field_type_5_is_host(
      meta_table_io_class_meta_init_bits_desc_state_field_type_5_is_host),
    .io_class_meta_init_bits_desc_state_field_type_6_is_repeated(
      meta_table_io_class_meta_init_bits_desc_state_field_type_6_is_repeated),
    .io_class_meta_init_bits_desc_state_field_type_6_field_type(
      meta_table_io_class_meta_init_bits_desc_state_field_type_6_field_type),
    .io_class_meta_init_bits_desc_state_field_type_6_sub_class_id(
      meta_table_io_class_meta_init_bits_desc_state_field_type_6_sub_class_id),
    .io_class_meta_init_bits_desc_state_field_type_6_is_host(
      meta_table_io_class_meta_init_bits_desc_state_field_type_6_is_host),
    .io_class_meta_init_bits_desc_state_field_type_7_is_repeated(
      meta_table_io_class_meta_init_bits_desc_state_field_type_7_is_repeated),
    .io_class_meta_init_bits_desc_state_field_type_7_field_type(
      meta_table_io_class_meta_init_bits_desc_state_field_type_7_field_type),
    .io_class_meta_init_bits_desc_state_field_type_7_sub_class_id(
      meta_table_io_class_meta_init_bits_desc_state_field_type_7_sub_class_id),
    .io_class_meta_init_bits_desc_state_field_type_7_is_host(
      meta_table_io_class_meta_init_bits_desc_state_field_type_7_is_host),
    .io_class_meta_init_bits_desc_state_field_type_8_is_repeated(
      meta_table_io_class_meta_init_bits_desc_state_field_type_8_is_repeated),
    .io_class_meta_init_bits_desc_state_field_type_8_field_type(
      meta_table_io_class_meta_init_bits_desc_state_field_type_8_field_type),
    .io_class_meta_init_bits_desc_state_field_type_8_sub_class_id(
      meta_table_io_class_meta_init_bits_desc_state_field_type_8_sub_class_id),
    .io_class_meta_init_bits_desc_state_field_type_8_is_host(
      meta_table_io_class_meta_init_bits_desc_state_field_type_8_is_host),
    .io_class_meta_init_bits_desc_state_field_type_9_is_repeated(
      meta_table_io_class_meta_init_bits_desc_state_field_type_9_is_repeated),
    .io_class_meta_init_bits_desc_state_field_type_9_field_type(
      meta_table_io_class_meta_init_bits_desc_state_field_type_9_field_type),
    .io_class_meta_init_bits_desc_state_field_type_9_sub_class_id(
      meta_table_io_class_meta_init_bits_desc_state_field_type_9_sub_class_id),
    .io_class_meta_init_bits_desc_state_field_type_9_is_host(
      meta_table_io_class_meta_init_bits_desc_state_field_type_9_is_host),
    .io_class_meta_init_bits_desc_state_field_type_10_is_repeated(
      meta_table_io_class_meta_init_bits_desc_state_field_type_10_is_repeated),
    .io_class_meta_init_bits_desc_state_field_type_10_field_type(
      meta_table_io_class_meta_init_bits_desc_state_field_type_10_field_type),
    .io_class_meta_init_bits_desc_state_field_type_10_sub_class_id(
      meta_table_io_class_meta_init_bits_desc_state_field_type_10_sub_class_id),
    .io_class_meta_init_bits_desc_state_field_type_10_is_host(
      meta_table_io_class_meta_init_bits_desc_state_field_type_10_is_host),
    .io_class_meta_init_bits_desc_state_field_type_11_is_repeated(
      meta_table_io_class_meta_init_bits_desc_state_field_type_11_is_repeated),
    .io_class_meta_init_bits_desc_state_field_type_11_field_type(
      meta_table_io_class_meta_init_bits_desc_state_field_type_11_field_type),
    .io_class_meta_init_bits_desc_state_field_type_11_sub_class_id(
      meta_table_io_class_meta_init_bits_desc_state_field_type_11_sub_class_id),
    .io_class_meta_init_bits_desc_state_field_type_11_is_host(
      meta_table_io_class_meta_init_bits_desc_state_field_type_11_is_host),
    .io_class_meta_init_bits_desc_state_field_type_12_is_repeated(
      meta_table_io_class_meta_init_bits_desc_state_field_type_12_is_repeated),
    .io_class_meta_init_bits_desc_state_field_type_12_field_type(
      meta_table_io_class_meta_init_bits_desc_state_field_type_12_field_type),
    .io_class_meta_init_bits_desc_state_field_type_12_sub_class_id(
      meta_table_io_class_meta_init_bits_desc_state_field_type_12_sub_class_id),
    .io_class_meta_init_bits_desc_state_field_type_12_is_host(
      meta_table_io_class_meta_init_bits_desc_state_field_type_12_is_host),
    .io_class_meta_init_bits_desc_state_field_type_13_is_repeated(
      meta_table_io_class_meta_init_bits_desc_state_field_type_13_is_repeated),
    .io_class_meta_init_bits_desc_state_field_type_13_field_type(
      meta_table_io_class_meta_init_bits_desc_state_field_type_13_field_type),
    .io_class_meta_init_bits_desc_state_field_type_13_sub_class_id(
      meta_table_io_class_meta_init_bits_desc_state_field_type_13_sub_class_id),
    .io_class_meta_init_bits_desc_state_field_type_13_is_host(
      meta_table_io_class_meta_init_bits_desc_state_field_type_13_is_host),
    .io_class_meta_init_bits_desc_state_field_type_14_is_repeated(
      meta_table_io_class_meta_init_bits_desc_state_field_type_14_is_repeated),
    .io_class_meta_init_bits_desc_state_field_type_14_field_type(
      meta_table_io_class_meta_init_bits_desc_state_field_type_14_field_type),
    .io_class_meta_init_bits_desc_state_field_type_14_sub_class_id(
      meta_table_io_class_meta_init_bits_desc_state_field_type_14_sub_class_id),
    .io_class_meta_init_bits_desc_state_field_type_14_is_host(
      meta_table_io_class_meta_init_bits_desc_state_field_type_14_is_host),
    .io_class_meta_init_bits_desc_state_field_type_15_is_repeated(
      meta_table_io_class_meta_init_bits_desc_state_field_type_15_is_repeated),
    .io_class_meta_init_bits_desc_state_field_type_15_field_type(
      meta_table_io_class_meta_init_bits_desc_state_field_type_15_field_type),
    .io_class_meta_init_bits_desc_state_field_type_15_sub_class_id(
      meta_table_io_class_meta_init_bits_desc_state_field_type_15_sub_class_id),
    .io_class_meta_init_bits_desc_state_field_type_15_is_host(
      meta_table_io_class_meta_init_bits_desc_state_field_type_15_is_host),
    .io_class_meta_init_bits_desc_state_field_type_16_is_repeated(
      meta_table_io_class_meta_init_bits_desc_state_field_type_16_is_repeated),
    .io_class_meta_init_bits_desc_state_field_type_16_field_type(
      meta_table_io_class_meta_init_bits_desc_state_field_type_16_field_type),
    .io_class_meta_init_bits_desc_state_field_type_16_sub_class_id(
      meta_table_io_class_meta_init_bits_desc_state_field_type_16_sub_class_id),
    .io_class_meta_init_bits_desc_state_field_type_16_is_host(
      meta_table_io_class_meta_init_bits_desc_state_field_type_16_is_host),
    .io_class_meta_init_bits_desc_state_field_type_17_is_repeated(
      meta_table_io_class_meta_init_bits_desc_state_field_type_17_is_repeated),
    .io_class_meta_init_bits_desc_state_field_type_17_field_type(
      meta_table_io_class_meta_init_bits_desc_state_field_type_17_field_type),
    .io_class_meta_init_bits_desc_state_field_type_17_sub_class_id(
      meta_table_io_class_meta_init_bits_desc_state_field_type_17_sub_class_id),
    .io_class_meta_init_bits_desc_state_field_type_17_is_host(
      meta_table_io_class_meta_init_bits_desc_state_field_type_17_is_host),
    .io_class_meta_init_bits_desc_state_field_type_18_is_repeated(
      meta_table_io_class_meta_init_bits_desc_state_field_type_18_is_repeated),
    .io_class_meta_init_bits_desc_state_field_type_18_field_type(
      meta_table_io_class_meta_init_bits_desc_state_field_type_18_field_type),
    .io_class_meta_init_bits_desc_state_field_type_18_sub_class_id(
      meta_table_io_class_meta_init_bits_desc_state_field_type_18_sub_class_id),
    .io_class_meta_init_bits_desc_state_field_type_18_is_host(
      meta_table_io_class_meta_init_bits_desc_state_field_type_18_is_host),
    .io_class_meta_init_bits_desc_state_field_type_19_is_repeated(
      meta_table_io_class_meta_init_bits_desc_state_field_type_19_is_repeated),
    .io_class_meta_init_bits_desc_state_field_type_19_field_type(
      meta_table_io_class_meta_init_bits_desc_state_field_type_19_field_type),
    .io_class_meta_init_bits_desc_state_field_type_19_sub_class_id(
      meta_table_io_class_meta_init_bits_desc_state_field_type_19_sub_class_id),
    .io_class_meta_init_bits_desc_state_field_type_19_is_host(
      meta_table_io_class_meta_init_bits_desc_state_field_type_19_is_host),
    .io_class_meta_init_bits_desc_state_field_type_20_is_repeated(
      meta_table_io_class_meta_init_bits_desc_state_field_type_20_is_repeated),
    .io_class_meta_init_bits_desc_state_field_type_20_field_type(
      meta_table_io_class_meta_init_bits_desc_state_field_type_20_field_type),
    .io_class_meta_init_bits_desc_state_field_type_20_sub_class_id(
      meta_table_io_class_meta_init_bits_desc_state_field_type_20_sub_class_id),
    .io_class_meta_init_bits_desc_state_field_type_20_is_host(
      meta_table_io_class_meta_init_bits_desc_state_field_type_20_is_host),
    .io_class_meta_init_bits_desc_state_field_type_21_is_repeated(
      meta_table_io_class_meta_init_bits_desc_state_field_type_21_is_repeated),
    .io_class_meta_init_bits_desc_state_field_type_21_field_type(
      meta_table_io_class_meta_init_bits_desc_state_field_type_21_field_type),
    .io_class_meta_init_bits_desc_state_field_type_21_sub_class_id(
      meta_table_io_class_meta_init_bits_desc_state_field_type_21_sub_class_id),
    .io_class_meta_init_bits_desc_state_field_type_21_is_host(
      meta_table_io_class_meta_init_bits_desc_state_field_type_21_is_host),
    .io_class_meta_init_bits_desc_state_field_type_22_is_repeated(
      meta_table_io_class_meta_init_bits_desc_state_field_type_22_is_repeated),
    .io_class_meta_init_bits_desc_state_field_type_22_field_type(
      meta_table_io_class_meta_init_bits_desc_state_field_type_22_field_type),
    .io_class_meta_init_bits_desc_state_field_type_22_sub_class_id(
      meta_table_io_class_meta_init_bits_desc_state_field_type_22_sub_class_id),
    .io_class_meta_init_bits_desc_state_field_type_22_is_host(
      meta_table_io_class_meta_init_bits_desc_state_field_type_22_is_host),
    .io_class_meta_init_bits_desc_state_field_type_23_is_repeated(
      meta_table_io_class_meta_init_bits_desc_state_field_type_23_is_repeated),
    .io_class_meta_init_bits_desc_state_field_type_23_field_type(
      meta_table_io_class_meta_init_bits_desc_state_field_type_23_field_type),
    .io_class_meta_init_bits_desc_state_field_type_23_sub_class_id(
      meta_table_io_class_meta_init_bits_desc_state_field_type_23_sub_class_id),
    .io_class_meta_init_bits_desc_state_field_type_23_is_host(
      meta_table_io_class_meta_init_bits_desc_state_field_type_23_is_host),
    .io_class_meta_init_bits_desc_state_field_type_24_is_repeated(
      meta_table_io_class_meta_init_bits_desc_state_field_type_24_is_repeated),
    .io_class_meta_init_bits_desc_state_field_type_24_field_type(
      meta_table_io_class_meta_init_bits_desc_state_field_type_24_field_type),
    .io_class_meta_init_bits_desc_state_field_type_24_sub_class_id(
      meta_table_io_class_meta_init_bits_desc_state_field_type_24_sub_class_id),
    .io_class_meta_init_bits_desc_state_field_type_24_is_host(
      meta_table_io_class_meta_init_bits_desc_state_field_type_24_is_host),
    .io_class_meta_init_bits_desc_state_field_type_25_is_repeated(
      meta_table_io_class_meta_init_bits_desc_state_field_type_25_is_repeated),
    .io_class_meta_init_bits_desc_state_field_type_25_field_type(
      meta_table_io_class_meta_init_bits_desc_state_field_type_25_field_type),
    .io_class_meta_init_bits_desc_state_field_type_25_sub_class_id(
      meta_table_io_class_meta_init_bits_desc_state_field_type_25_sub_class_id),
    .io_class_meta_init_bits_desc_state_field_type_25_is_host(
      meta_table_io_class_meta_init_bits_desc_state_field_type_25_is_host),
    .io_class_meta_init_bits_desc_state_field_type_26_is_repeated(
      meta_table_io_class_meta_init_bits_desc_state_field_type_26_is_repeated),
    .io_class_meta_init_bits_desc_state_field_type_26_field_type(
      meta_table_io_class_meta_init_bits_desc_state_field_type_26_field_type),
    .io_class_meta_init_bits_desc_state_field_type_26_sub_class_id(
      meta_table_io_class_meta_init_bits_desc_state_field_type_26_sub_class_id),
    .io_class_meta_init_bits_desc_state_field_type_26_is_host(
      meta_table_io_class_meta_init_bits_desc_state_field_type_26_is_host),
    .io_class_meta_init_bits_desc_state_field_type_27_is_repeated(
      meta_table_io_class_meta_init_bits_desc_state_field_type_27_is_repeated),
    .io_class_meta_init_bits_desc_state_field_type_27_field_type(
      meta_table_io_class_meta_init_bits_desc_state_field_type_27_field_type),
    .io_class_meta_init_bits_desc_state_field_type_27_sub_class_id(
      meta_table_io_class_meta_init_bits_desc_state_field_type_27_sub_class_id),
    .io_class_meta_init_bits_desc_state_field_type_27_is_host(
      meta_table_io_class_meta_init_bits_desc_state_field_type_27_is_host),
    .io_class_meta_init_bits_desc_state_field_type_28_is_repeated(
      meta_table_io_class_meta_init_bits_desc_state_field_type_28_is_repeated),
    .io_class_meta_init_bits_desc_state_field_type_28_field_type(
      meta_table_io_class_meta_init_bits_desc_state_field_type_28_field_type),
    .io_class_meta_init_bits_desc_state_field_type_28_sub_class_id(
      meta_table_io_class_meta_init_bits_desc_state_field_type_28_sub_class_id),
    .io_class_meta_init_bits_desc_state_field_type_28_is_host(
      meta_table_io_class_meta_init_bits_desc_state_field_type_28_is_host),
    .io_class_meta_init_bits_desc_state_field_type_29_is_repeated(
      meta_table_io_class_meta_init_bits_desc_state_field_type_29_is_repeated),
    .io_class_meta_init_bits_desc_state_field_type_29_field_type(
      meta_table_io_class_meta_init_bits_desc_state_field_type_29_field_type),
    .io_class_meta_init_bits_desc_state_field_type_29_sub_class_id(
      meta_table_io_class_meta_init_bits_desc_state_field_type_29_sub_class_id),
    .io_class_meta_init_bits_desc_state_field_type_29_is_host(
      meta_table_io_class_meta_init_bits_desc_state_field_type_29_is_host),
    .io_class_meta_init_bits_desc_state_field_type_30_is_repeated(
      meta_table_io_class_meta_init_bits_desc_state_field_type_30_is_repeated),
    .io_class_meta_init_bits_desc_state_field_type_30_field_type(
      meta_table_io_class_meta_init_bits_desc_state_field_type_30_field_type),
    .io_class_meta_init_bits_desc_state_field_type_30_sub_class_id(
      meta_table_io_class_meta_init_bits_desc_state_field_type_30_sub_class_id),
    .io_class_meta_init_bits_desc_state_field_type_30_is_host(
      meta_table_io_class_meta_init_bits_desc_state_field_type_30_is_host),
    .io_class_meta_init_bits_desc_state_field_type_31_is_repeated(
      meta_table_io_class_meta_init_bits_desc_state_field_type_31_is_repeated),
    .io_class_meta_init_bits_desc_state_field_type_31_field_type(
      meta_table_io_class_meta_init_bits_desc_state_field_type_31_field_type),
    .io_class_meta_init_bits_desc_state_field_type_31_sub_class_id(
      meta_table_io_class_meta_init_bits_desc_state_field_type_31_sub_class_id),
    .io_class_meta_init_bits_desc_state_field_type_31_is_host(
      meta_table_io_class_meta_init_bits_desc_state_field_type_31_is_host),
    .io_class_meta_init_bits_desc_state_field_type_32_is_repeated(
      meta_table_io_class_meta_init_bits_desc_state_field_type_32_is_repeated),
    .io_class_meta_init_bits_desc_state_field_type_32_field_type(
      meta_table_io_class_meta_init_bits_desc_state_field_type_32_field_type),
    .io_class_meta_init_bits_desc_state_field_type_32_sub_class_id(
      meta_table_io_class_meta_init_bits_desc_state_field_type_32_sub_class_id),
    .io_class_meta_init_bits_desc_state_field_type_32_is_host(
      meta_table_io_class_meta_init_bits_desc_state_field_type_32_is_host),
    .io_s_class_meta_req_ready(meta_table_io_s_class_meta_req_ready),
    .io_s_class_meta_req_valid(meta_table_io_s_class_meta_req_valid),
    .io_s_class_meta_req_bits_class_id(meta_table_io_s_class_meta_req_bits_class_id),
    .io_s_class_meta_rsp_valid(meta_table_io_s_class_meta_rsp_valid),
    .io_s_class_meta_rsp_bits_class_meta_max_field_num(meta_table_io_s_class_meta_rsp_bits_class_meta_max_field_num),
    .io_s_class_meta_rsp_bits_class_meta_field_type_0_is_repeated(
      meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_0_is_repeated),
    .io_s_class_meta_rsp_bits_class_meta_field_type_0_field_type(
      meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_0_field_type),
    .io_s_class_meta_rsp_bits_class_meta_field_type_0_sub_class_id(
      meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_0_sub_class_id),
    .io_s_class_meta_rsp_bits_class_meta_field_type_1_is_repeated(
      meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_1_is_repeated),
    .io_s_class_meta_rsp_bits_class_meta_field_type_1_field_type(
      meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_1_field_type),
    .io_s_class_meta_rsp_bits_class_meta_field_type_1_sub_class_id(
      meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_1_sub_class_id),
    .io_s_class_meta_rsp_bits_class_meta_field_type_2_is_repeated(
      meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_2_is_repeated),
    .io_s_class_meta_rsp_bits_class_meta_field_type_2_field_type(
      meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_2_field_type),
    .io_s_class_meta_rsp_bits_class_meta_field_type_2_sub_class_id(
      meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_2_sub_class_id),
    .io_s_class_meta_rsp_bits_class_meta_field_type_3_is_repeated(
      meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_3_is_repeated),
    .io_s_class_meta_rsp_bits_class_meta_field_type_3_field_type(
      meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_3_field_type),
    .io_s_class_meta_rsp_bits_class_meta_field_type_3_sub_class_id(
      meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_3_sub_class_id),
    .io_s_class_meta_rsp_bits_class_meta_field_type_4_is_repeated(
      meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_4_is_repeated),
    .io_s_class_meta_rsp_bits_class_meta_field_type_4_field_type(
      meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_4_field_type),
    .io_s_class_meta_rsp_bits_class_meta_field_type_4_sub_class_id(
      meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_4_sub_class_id),
    .io_s_class_meta_rsp_bits_class_meta_field_type_5_is_repeated(
      meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_5_is_repeated),
    .io_s_class_meta_rsp_bits_class_meta_field_type_5_field_type(
      meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_5_field_type),
    .io_s_class_meta_rsp_bits_class_meta_field_type_5_sub_class_id(
      meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_5_sub_class_id),
    .io_s_class_meta_rsp_bits_class_meta_field_type_6_is_repeated(
      meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_6_is_repeated),
    .io_s_class_meta_rsp_bits_class_meta_field_type_6_field_type(
      meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_6_field_type),
    .io_s_class_meta_rsp_bits_class_meta_field_type_6_sub_class_id(
      meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_6_sub_class_id),
    .io_s_class_meta_rsp_bits_class_meta_field_type_7_is_repeated(
      meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_7_is_repeated),
    .io_s_class_meta_rsp_bits_class_meta_field_type_7_field_type(
      meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_7_field_type),
    .io_s_class_meta_rsp_bits_class_meta_field_type_7_sub_class_id(
      meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_7_sub_class_id),
    .io_s_class_meta_rsp_bits_class_meta_field_type_8_is_repeated(
      meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_8_is_repeated),
    .io_s_class_meta_rsp_bits_class_meta_field_type_8_field_type(
      meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_8_field_type),
    .io_s_class_meta_rsp_bits_class_meta_field_type_8_sub_class_id(
      meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_8_sub_class_id),
    .io_s_class_meta_rsp_bits_class_meta_field_type_9_is_repeated(
      meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_9_is_repeated),
    .io_s_class_meta_rsp_bits_class_meta_field_type_9_field_type(
      meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_9_field_type),
    .io_s_class_meta_rsp_bits_class_meta_field_type_9_sub_class_id(
      meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_9_sub_class_id),
    .io_s_class_meta_rsp_bits_class_meta_field_type_10_is_repeated(
      meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_10_is_repeated),
    .io_s_class_meta_rsp_bits_class_meta_field_type_10_field_type(
      meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_10_field_type),
    .io_s_class_meta_rsp_bits_class_meta_field_type_10_sub_class_id(
      meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_10_sub_class_id),
    .io_s_class_meta_rsp_bits_class_meta_field_type_11_is_repeated(
      meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_11_is_repeated),
    .io_s_class_meta_rsp_bits_class_meta_field_type_11_field_type(
      meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_11_field_type),
    .io_s_class_meta_rsp_bits_class_meta_field_type_11_sub_class_id(
      meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_11_sub_class_id),
    .io_s_class_meta_rsp_bits_class_meta_field_type_12_is_repeated(
      meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_12_is_repeated),
    .io_s_class_meta_rsp_bits_class_meta_field_type_12_field_type(
      meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_12_field_type),
    .io_s_class_meta_rsp_bits_class_meta_field_type_12_sub_class_id(
      meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_12_sub_class_id),
    .io_s_class_meta_rsp_bits_class_meta_field_type_13_is_repeated(
      meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_13_is_repeated),
    .io_s_class_meta_rsp_bits_class_meta_field_type_13_field_type(
      meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_13_field_type),
    .io_s_class_meta_rsp_bits_class_meta_field_type_13_sub_class_id(
      meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_13_sub_class_id),
    .io_s_class_meta_rsp_bits_class_meta_field_type_14_is_repeated(
      meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_14_is_repeated),
    .io_s_class_meta_rsp_bits_class_meta_field_type_14_field_type(
      meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_14_field_type),
    .io_s_class_meta_rsp_bits_class_meta_field_type_14_sub_class_id(
      meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_14_sub_class_id),
    .io_s_class_meta_rsp_bits_class_meta_field_type_15_is_repeated(
      meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_15_is_repeated),
    .io_s_class_meta_rsp_bits_class_meta_field_type_15_field_type(
      meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_15_field_type),
    .io_s_class_meta_rsp_bits_class_meta_field_type_15_sub_class_id(
      meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_15_sub_class_id),
    .io_s_class_meta_rsp_bits_class_meta_field_type_16_is_repeated(
      meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_16_is_repeated),
    .io_s_class_meta_rsp_bits_class_meta_field_type_16_field_type(
      meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_16_field_type),
    .io_s_class_meta_rsp_bits_class_meta_field_type_16_sub_class_id(
      meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_16_sub_class_id),
    .io_s_class_meta_rsp_bits_class_meta_field_type_17_is_repeated(
      meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_17_is_repeated),
    .io_s_class_meta_rsp_bits_class_meta_field_type_17_field_type(
      meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_17_field_type),
    .io_s_class_meta_rsp_bits_class_meta_field_type_17_sub_class_id(
      meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_17_sub_class_id),
    .io_s_class_meta_rsp_bits_class_meta_field_type_18_is_repeated(
      meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_18_is_repeated),
    .io_s_class_meta_rsp_bits_class_meta_field_type_18_field_type(
      meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_18_field_type),
    .io_s_class_meta_rsp_bits_class_meta_field_type_18_sub_class_id(
      meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_18_sub_class_id),
    .io_s_class_meta_rsp_bits_class_meta_field_type_19_is_repeated(
      meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_19_is_repeated),
    .io_s_class_meta_rsp_bits_class_meta_field_type_19_field_type(
      meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_19_field_type),
    .io_s_class_meta_rsp_bits_class_meta_field_type_19_sub_class_id(
      meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_19_sub_class_id),
    .io_s_class_meta_rsp_bits_class_meta_field_type_20_is_repeated(
      meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_20_is_repeated),
    .io_s_class_meta_rsp_bits_class_meta_field_type_20_field_type(
      meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_20_field_type),
    .io_s_class_meta_rsp_bits_class_meta_field_type_20_sub_class_id(
      meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_20_sub_class_id),
    .io_s_class_meta_rsp_bits_class_meta_field_type_21_is_repeated(
      meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_21_is_repeated),
    .io_s_class_meta_rsp_bits_class_meta_field_type_21_field_type(
      meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_21_field_type),
    .io_s_class_meta_rsp_bits_class_meta_field_type_21_sub_class_id(
      meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_21_sub_class_id),
    .io_s_class_meta_rsp_bits_class_meta_field_type_22_is_repeated(
      meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_22_is_repeated),
    .io_s_class_meta_rsp_bits_class_meta_field_type_22_field_type(
      meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_22_field_type),
    .io_s_class_meta_rsp_bits_class_meta_field_type_22_sub_class_id(
      meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_22_sub_class_id),
    .io_s_class_meta_rsp_bits_class_meta_field_type_23_is_repeated(
      meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_23_is_repeated),
    .io_s_class_meta_rsp_bits_class_meta_field_type_23_field_type(
      meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_23_field_type),
    .io_s_class_meta_rsp_bits_class_meta_field_type_23_sub_class_id(
      meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_23_sub_class_id),
    .io_s_class_meta_rsp_bits_class_meta_field_type_24_is_repeated(
      meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_24_is_repeated),
    .io_s_class_meta_rsp_bits_class_meta_field_type_24_field_type(
      meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_24_field_type),
    .io_s_class_meta_rsp_bits_class_meta_field_type_24_sub_class_id(
      meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_24_sub_class_id),
    .io_s_class_meta_rsp_bits_class_meta_field_type_25_is_repeated(
      meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_25_is_repeated),
    .io_s_class_meta_rsp_bits_class_meta_field_type_25_field_type(
      meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_25_field_type),
    .io_s_class_meta_rsp_bits_class_meta_field_type_25_sub_class_id(
      meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_25_sub_class_id),
    .io_s_class_meta_rsp_bits_class_meta_field_type_26_is_repeated(
      meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_26_is_repeated),
    .io_s_class_meta_rsp_bits_class_meta_field_type_26_field_type(
      meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_26_field_type),
    .io_s_class_meta_rsp_bits_class_meta_field_type_26_sub_class_id(
      meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_26_sub_class_id),
    .io_s_class_meta_rsp_bits_class_meta_field_type_27_is_repeated(
      meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_27_is_repeated),
    .io_s_class_meta_rsp_bits_class_meta_field_type_27_field_type(
      meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_27_field_type),
    .io_s_class_meta_rsp_bits_class_meta_field_type_27_sub_class_id(
      meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_27_sub_class_id),
    .io_s_class_meta_rsp_bits_class_meta_field_type_28_is_repeated(
      meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_28_is_repeated),
    .io_s_class_meta_rsp_bits_class_meta_field_type_28_field_type(
      meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_28_field_type),
    .io_s_class_meta_rsp_bits_class_meta_field_type_28_sub_class_id(
      meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_28_sub_class_id),
    .io_s_class_meta_rsp_bits_class_meta_field_type_29_is_repeated(
      meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_29_is_repeated),
    .io_s_class_meta_rsp_bits_class_meta_field_type_29_field_type(
      meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_29_field_type),
    .io_s_class_meta_rsp_bits_class_meta_field_type_29_sub_class_id(
      meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_29_sub_class_id),
    .io_s_class_meta_rsp_bits_class_meta_field_type_30_is_repeated(
      meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_30_is_repeated),
    .io_s_class_meta_rsp_bits_class_meta_field_type_30_field_type(
      meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_30_field_type),
    .io_s_class_meta_rsp_bits_class_meta_field_type_30_sub_class_id(
      meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_30_sub_class_id),
    .io_s_class_meta_rsp_bits_class_meta_field_type_31_is_repeated(
      meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_31_is_repeated),
    .io_s_class_meta_rsp_bits_class_meta_field_type_31_field_type(
      meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_31_field_type),
    .io_s_class_meta_rsp_bits_class_meta_field_type_31_sub_class_id(
      meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_31_sub_class_id),
    .io_s_class_meta_rsp_bits_class_meta_field_type_32_is_repeated(
      meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_32_is_repeated),
    .io_s_class_meta_rsp_bits_class_meta_field_type_32_field_type(
      meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_32_field_type),
    .io_s_class_meta_rsp_bits_class_meta_field_type_32_sub_class_id(
      meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_32_sub_class_id),
    .counter_5(meta_table_counter_5)
  );
  Control control ( // @[FpgaCloudSerHw.scala 108:29]
    .clock(control_clock),
    .reset(control_reset),
    .io_axi_aw_ready(control_io_axi_aw_ready),
    .io_axi_aw_valid(control_io_axi_aw_valid),
    .io_axi_aw_bits_addr(control_io_axi_aw_bits_addr),
    .io_axi_w_ready(control_io_axi_w_ready),
    .io_axi_w_valid(control_io_axi_w_valid),
    .io_axi_w_bits_data(control_io_axi_w_bits_data),
    .io_axi_r_ready(control_io_axi_r_ready),
    .io_axi_r_valid(control_io_axi_r_valid),
    .io_axi_r_bits_data(control_io_axi_r_bits_data),
    .io_metadata_init_valid(control_io_metadata_init_valid),
    .io_metadata_init_bits_class_id(control_io_metadata_init_bits_class_id),
    .io_metadata_init_bits_desc_state_class_length(control_io_metadata_init_bits_desc_state_class_length),
    .io_metadata_init_bits_desc_state_max_field_num(control_io_metadata_init_bits_desc_state_max_field_num),
    .io_metadata_init_bits_desc_state_field_type_0_is_repeated(
      control_io_metadata_init_bits_desc_state_field_type_0_is_repeated),
    .io_metadata_init_bits_desc_state_field_type_0_field_type(
      control_io_metadata_init_bits_desc_state_field_type_0_field_type),
    .io_metadata_init_bits_desc_state_field_type_0_sub_class_id(
      control_io_metadata_init_bits_desc_state_field_type_0_sub_class_id),
    .io_metadata_init_bits_desc_state_field_type_0_is_host(control_io_metadata_init_bits_desc_state_field_type_0_is_host
      ),
    .io_metadata_init_bits_desc_state_field_type_1_is_repeated(
      control_io_metadata_init_bits_desc_state_field_type_1_is_repeated),
    .io_metadata_init_bits_desc_state_field_type_1_field_type(
      control_io_metadata_init_bits_desc_state_field_type_1_field_type),
    .io_metadata_init_bits_desc_state_field_type_1_sub_class_id(
      control_io_metadata_init_bits_desc_state_field_type_1_sub_class_id),
    .io_metadata_init_bits_desc_state_field_type_1_is_host(control_io_metadata_init_bits_desc_state_field_type_1_is_host
      ),
    .io_metadata_init_bits_desc_state_field_type_2_is_repeated(
      control_io_metadata_init_bits_desc_state_field_type_2_is_repeated),
    .io_metadata_init_bits_desc_state_field_type_2_field_type(
      control_io_metadata_init_bits_desc_state_field_type_2_field_type),
    .io_metadata_init_bits_desc_state_field_type_2_sub_class_id(
      control_io_metadata_init_bits_desc_state_field_type_2_sub_class_id),
    .io_metadata_init_bits_desc_state_field_type_2_is_host(control_io_metadata_init_bits_desc_state_field_type_2_is_host
      ),
    .io_metadata_init_bits_desc_state_field_type_3_is_repeated(
      control_io_metadata_init_bits_desc_state_field_type_3_is_repeated),
    .io_metadata_init_bits_desc_state_field_type_3_field_type(
      control_io_metadata_init_bits_desc_state_field_type_3_field_type),
    .io_metadata_init_bits_desc_state_field_type_3_sub_class_id(
      control_io_metadata_init_bits_desc_state_field_type_3_sub_class_id),
    .io_metadata_init_bits_desc_state_field_type_3_is_host(control_io_metadata_init_bits_desc_state_field_type_3_is_host
      ),
    .io_metadata_init_bits_desc_state_field_type_4_is_repeated(
      control_io_metadata_init_bits_desc_state_field_type_4_is_repeated),
    .io_metadata_init_bits_desc_state_field_type_4_field_type(
      control_io_metadata_init_bits_desc_state_field_type_4_field_type),
    .io_metadata_init_bits_desc_state_field_type_4_sub_class_id(
      control_io_metadata_init_bits_desc_state_field_type_4_sub_class_id),
    .io_metadata_init_bits_desc_state_field_type_4_is_host(control_io_metadata_init_bits_desc_state_field_type_4_is_host
      ),
    .io_metadata_init_bits_desc_state_field_type_5_is_repeated(
      control_io_metadata_init_bits_desc_state_field_type_5_is_repeated),
    .io_metadata_init_bits_desc_state_field_type_5_field_type(
      control_io_metadata_init_bits_desc_state_field_type_5_field_type),
    .io_metadata_init_bits_desc_state_field_type_5_sub_class_id(
      control_io_metadata_init_bits_desc_state_field_type_5_sub_class_id),
    .io_metadata_init_bits_desc_state_field_type_5_is_host(control_io_metadata_init_bits_desc_state_field_type_5_is_host
      ),
    .io_metadata_init_bits_desc_state_field_type_6_is_repeated(
      control_io_metadata_init_bits_desc_state_field_type_6_is_repeated),
    .io_metadata_init_bits_desc_state_field_type_6_field_type(
      control_io_metadata_init_bits_desc_state_field_type_6_field_type),
    .io_metadata_init_bits_desc_state_field_type_6_sub_class_id(
      control_io_metadata_init_bits_desc_state_field_type_6_sub_class_id),
    .io_metadata_init_bits_desc_state_field_type_6_is_host(control_io_metadata_init_bits_desc_state_field_type_6_is_host
      ),
    .io_metadata_init_bits_desc_state_field_type_7_is_repeated(
      control_io_metadata_init_bits_desc_state_field_type_7_is_repeated),
    .io_metadata_init_bits_desc_state_field_type_7_field_type(
      control_io_metadata_init_bits_desc_state_field_type_7_field_type),
    .io_metadata_init_bits_desc_state_field_type_7_sub_class_id(
      control_io_metadata_init_bits_desc_state_field_type_7_sub_class_id),
    .io_metadata_init_bits_desc_state_field_type_7_is_host(control_io_metadata_init_bits_desc_state_field_type_7_is_host
      ),
    .io_metadata_init_bits_desc_state_field_type_8_is_repeated(
      control_io_metadata_init_bits_desc_state_field_type_8_is_repeated),
    .io_metadata_init_bits_desc_state_field_type_8_field_type(
      control_io_metadata_init_bits_desc_state_field_type_8_field_type),
    .io_metadata_init_bits_desc_state_field_type_8_sub_class_id(
      control_io_metadata_init_bits_desc_state_field_type_8_sub_class_id),
    .io_metadata_init_bits_desc_state_field_type_8_is_host(control_io_metadata_init_bits_desc_state_field_type_8_is_host
      ),
    .io_metadata_init_bits_desc_state_field_type_9_is_repeated(
      control_io_metadata_init_bits_desc_state_field_type_9_is_repeated),
    .io_metadata_init_bits_desc_state_field_type_9_field_type(
      control_io_metadata_init_bits_desc_state_field_type_9_field_type),
    .io_metadata_init_bits_desc_state_field_type_9_sub_class_id(
      control_io_metadata_init_bits_desc_state_field_type_9_sub_class_id),
    .io_metadata_init_bits_desc_state_field_type_9_is_host(control_io_metadata_init_bits_desc_state_field_type_9_is_host
      ),
    .io_metadata_init_bits_desc_state_field_type_10_is_repeated(
      control_io_metadata_init_bits_desc_state_field_type_10_is_repeated),
    .io_metadata_init_bits_desc_state_field_type_10_field_type(
      control_io_metadata_init_bits_desc_state_field_type_10_field_type),
    .io_metadata_init_bits_desc_state_field_type_10_sub_class_id(
      control_io_metadata_init_bits_desc_state_field_type_10_sub_class_id),
    .io_metadata_init_bits_desc_state_field_type_10_is_host(
      control_io_metadata_init_bits_desc_state_field_type_10_is_host),
    .io_metadata_init_bits_desc_state_field_type_11_is_repeated(
      control_io_metadata_init_bits_desc_state_field_type_11_is_repeated),
    .io_metadata_init_bits_desc_state_field_type_11_field_type(
      control_io_metadata_init_bits_desc_state_field_type_11_field_type),
    .io_metadata_init_bits_desc_state_field_type_11_sub_class_id(
      control_io_metadata_init_bits_desc_state_field_type_11_sub_class_id),
    .io_metadata_init_bits_desc_state_field_type_11_is_host(
      control_io_metadata_init_bits_desc_state_field_type_11_is_host),
    .io_metadata_init_bits_desc_state_field_type_12_is_repeated(
      control_io_metadata_init_bits_desc_state_field_type_12_is_repeated),
    .io_metadata_init_bits_desc_state_field_type_12_field_type(
      control_io_metadata_init_bits_desc_state_field_type_12_field_type),
    .io_metadata_init_bits_desc_state_field_type_12_sub_class_id(
      control_io_metadata_init_bits_desc_state_field_type_12_sub_class_id),
    .io_metadata_init_bits_desc_state_field_type_12_is_host(
      control_io_metadata_init_bits_desc_state_field_type_12_is_host),
    .io_metadata_init_bits_desc_state_field_type_13_is_repeated(
      control_io_metadata_init_bits_desc_state_field_type_13_is_repeated),
    .io_metadata_init_bits_desc_state_field_type_13_field_type(
      control_io_metadata_init_bits_desc_state_field_type_13_field_type),
    .io_metadata_init_bits_desc_state_field_type_13_sub_class_id(
      control_io_metadata_init_bits_desc_state_field_type_13_sub_class_id),
    .io_metadata_init_bits_desc_state_field_type_13_is_host(
      control_io_metadata_init_bits_desc_state_field_type_13_is_host),
    .io_metadata_init_bits_desc_state_field_type_14_is_repeated(
      control_io_metadata_init_bits_desc_state_field_type_14_is_repeated),
    .io_metadata_init_bits_desc_state_field_type_14_field_type(
      control_io_metadata_init_bits_desc_state_field_type_14_field_type),
    .io_metadata_init_bits_desc_state_field_type_14_sub_class_id(
      control_io_metadata_init_bits_desc_state_field_type_14_sub_class_id),
    .io_metadata_init_bits_desc_state_field_type_14_is_host(
      control_io_metadata_init_bits_desc_state_field_type_14_is_host),
    .io_metadata_init_bits_desc_state_field_type_15_is_repeated(
      control_io_metadata_init_bits_desc_state_field_type_15_is_repeated),
    .io_metadata_init_bits_desc_state_field_type_15_field_type(
      control_io_metadata_init_bits_desc_state_field_type_15_field_type),
    .io_metadata_init_bits_desc_state_field_type_15_sub_class_id(
      control_io_metadata_init_bits_desc_state_field_type_15_sub_class_id),
    .io_metadata_init_bits_desc_state_field_type_15_is_host(
      control_io_metadata_init_bits_desc_state_field_type_15_is_host),
    .io_metadata_init_bits_desc_state_field_type_16_is_repeated(
      control_io_metadata_init_bits_desc_state_field_type_16_is_repeated),
    .io_metadata_init_bits_desc_state_field_type_16_field_type(
      control_io_metadata_init_bits_desc_state_field_type_16_field_type),
    .io_metadata_init_bits_desc_state_field_type_16_sub_class_id(
      control_io_metadata_init_bits_desc_state_field_type_16_sub_class_id),
    .io_metadata_init_bits_desc_state_field_type_16_is_host(
      control_io_metadata_init_bits_desc_state_field_type_16_is_host),
    .io_metadata_init_bits_desc_state_field_type_17_is_repeated(
      control_io_metadata_init_bits_desc_state_field_type_17_is_repeated),
    .io_metadata_init_bits_desc_state_field_type_17_field_type(
      control_io_metadata_init_bits_desc_state_field_type_17_field_type),
    .io_metadata_init_bits_desc_state_field_type_17_sub_class_id(
      control_io_metadata_init_bits_desc_state_field_type_17_sub_class_id),
    .io_metadata_init_bits_desc_state_field_type_17_is_host(
      control_io_metadata_init_bits_desc_state_field_type_17_is_host),
    .io_metadata_init_bits_desc_state_field_type_18_is_repeated(
      control_io_metadata_init_bits_desc_state_field_type_18_is_repeated),
    .io_metadata_init_bits_desc_state_field_type_18_field_type(
      control_io_metadata_init_bits_desc_state_field_type_18_field_type),
    .io_metadata_init_bits_desc_state_field_type_18_sub_class_id(
      control_io_metadata_init_bits_desc_state_field_type_18_sub_class_id),
    .io_metadata_init_bits_desc_state_field_type_18_is_host(
      control_io_metadata_init_bits_desc_state_field_type_18_is_host),
    .io_metadata_init_bits_desc_state_field_type_19_is_repeated(
      control_io_metadata_init_bits_desc_state_field_type_19_is_repeated),
    .io_metadata_init_bits_desc_state_field_type_19_field_type(
      control_io_metadata_init_bits_desc_state_field_type_19_field_type),
    .io_metadata_init_bits_desc_state_field_type_19_sub_class_id(
      control_io_metadata_init_bits_desc_state_field_type_19_sub_class_id),
    .io_metadata_init_bits_desc_state_field_type_19_is_host(
      control_io_metadata_init_bits_desc_state_field_type_19_is_host),
    .io_metadata_init_bits_desc_state_field_type_20_is_repeated(
      control_io_metadata_init_bits_desc_state_field_type_20_is_repeated),
    .io_metadata_init_bits_desc_state_field_type_20_field_type(
      control_io_metadata_init_bits_desc_state_field_type_20_field_type),
    .io_metadata_init_bits_desc_state_field_type_20_sub_class_id(
      control_io_metadata_init_bits_desc_state_field_type_20_sub_class_id),
    .io_metadata_init_bits_desc_state_field_type_20_is_host(
      control_io_metadata_init_bits_desc_state_field_type_20_is_host),
    .io_metadata_init_bits_desc_state_field_type_21_is_repeated(
      control_io_metadata_init_bits_desc_state_field_type_21_is_repeated),
    .io_metadata_init_bits_desc_state_field_type_21_field_type(
      control_io_metadata_init_bits_desc_state_field_type_21_field_type),
    .io_metadata_init_bits_desc_state_field_type_21_sub_class_id(
      control_io_metadata_init_bits_desc_state_field_type_21_sub_class_id),
    .io_metadata_init_bits_desc_state_field_type_21_is_host(
      control_io_metadata_init_bits_desc_state_field_type_21_is_host),
    .io_metadata_init_bits_desc_state_field_type_22_is_repeated(
      control_io_metadata_init_bits_desc_state_field_type_22_is_repeated),
    .io_metadata_init_bits_desc_state_field_type_22_field_type(
      control_io_metadata_init_bits_desc_state_field_type_22_field_type),
    .io_metadata_init_bits_desc_state_field_type_22_sub_class_id(
      control_io_metadata_init_bits_desc_state_field_type_22_sub_class_id),
    .io_metadata_init_bits_desc_state_field_type_22_is_host(
      control_io_metadata_init_bits_desc_state_field_type_22_is_host),
    .io_metadata_init_bits_desc_state_field_type_23_is_repeated(
      control_io_metadata_init_bits_desc_state_field_type_23_is_repeated),
    .io_metadata_init_bits_desc_state_field_type_23_field_type(
      control_io_metadata_init_bits_desc_state_field_type_23_field_type),
    .io_metadata_init_bits_desc_state_field_type_23_sub_class_id(
      control_io_metadata_init_bits_desc_state_field_type_23_sub_class_id),
    .io_metadata_init_bits_desc_state_field_type_23_is_host(
      control_io_metadata_init_bits_desc_state_field_type_23_is_host),
    .io_metadata_init_bits_desc_state_field_type_24_is_repeated(
      control_io_metadata_init_bits_desc_state_field_type_24_is_repeated),
    .io_metadata_init_bits_desc_state_field_type_24_field_type(
      control_io_metadata_init_bits_desc_state_field_type_24_field_type),
    .io_metadata_init_bits_desc_state_field_type_24_sub_class_id(
      control_io_metadata_init_bits_desc_state_field_type_24_sub_class_id),
    .io_metadata_init_bits_desc_state_field_type_24_is_host(
      control_io_metadata_init_bits_desc_state_field_type_24_is_host),
    .io_metadata_init_bits_desc_state_field_type_25_is_repeated(
      control_io_metadata_init_bits_desc_state_field_type_25_is_repeated),
    .io_metadata_init_bits_desc_state_field_type_25_field_type(
      control_io_metadata_init_bits_desc_state_field_type_25_field_type),
    .io_metadata_init_bits_desc_state_field_type_25_sub_class_id(
      control_io_metadata_init_bits_desc_state_field_type_25_sub_class_id),
    .io_metadata_init_bits_desc_state_field_type_25_is_host(
      control_io_metadata_init_bits_desc_state_field_type_25_is_host),
    .io_metadata_init_bits_desc_state_field_type_26_is_repeated(
      control_io_metadata_init_bits_desc_state_field_type_26_is_repeated),
    .io_metadata_init_bits_desc_state_field_type_26_field_type(
      control_io_metadata_init_bits_desc_state_field_type_26_field_type),
    .io_metadata_init_bits_desc_state_field_type_26_sub_class_id(
      control_io_metadata_init_bits_desc_state_field_type_26_sub_class_id),
    .io_metadata_init_bits_desc_state_field_type_26_is_host(
      control_io_metadata_init_bits_desc_state_field_type_26_is_host),
    .io_metadata_init_bits_desc_state_field_type_27_is_repeated(
      control_io_metadata_init_bits_desc_state_field_type_27_is_repeated),
    .io_metadata_init_bits_desc_state_field_type_27_field_type(
      control_io_metadata_init_bits_desc_state_field_type_27_field_type),
    .io_metadata_init_bits_desc_state_field_type_27_sub_class_id(
      control_io_metadata_init_bits_desc_state_field_type_27_sub_class_id),
    .io_metadata_init_bits_desc_state_field_type_27_is_host(
      control_io_metadata_init_bits_desc_state_field_type_27_is_host),
    .io_metadata_init_bits_desc_state_field_type_28_is_repeated(
      control_io_metadata_init_bits_desc_state_field_type_28_is_repeated),
    .io_metadata_init_bits_desc_state_field_type_28_field_type(
      control_io_metadata_init_bits_desc_state_field_type_28_field_type),
    .io_metadata_init_bits_desc_state_field_type_28_sub_class_id(
      control_io_metadata_init_bits_desc_state_field_type_28_sub_class_id),
    .io_metadata_init_bits_desc_state_field_type_28_is_host(
      control_io_metadata_init_bits_desc_state_field_type_28_is_host),
    .io_metadata_init_bits_desc_state_field_type_29_is_repeated(
      control_io_metadata_init_bits_desc_state_field_type_29_is_repeated),
    .io_metadata_init_bits_desc_state_field_type_29_field_type(
      control_io_metadata_init_bits_desc_state_field_type_29_field_type),
    .io_metadata_init_bits_desc_state_field_type_29_sub_class_id(
      control_io_metadata_init_bits_desc_state_field_type_29_sub_class_id),
    .io_metadata_init_bits_desc_state_field_type_29_is_host(
      control_io_metadata_init_bits_desc_state_field_type_29_is_host),
    .io_metadata_init_bits_desc_state_field_type_30_is_repeated(
      control_io_metadata_init_bits_desc_state_field_type_30_is_repeated),
    .io_metadata_init_bits_desc_state_field_type_30_field_type(
      control_io_metadata_init_bits_desc_state_field_type_30_field_type),
    .io_metadata_init_bits_desc_state_field_type_30_sub_class_id(
      control_io_metadata_init_bits_desc_state_field_type_30_sub_class_id),
    .io_metadata_init_bits_desc_state_field_type_30_is_host(
      control_io_metadata_init_bits_desc_state_field_type_30_is_host),
    .io_metadata_init_bits_desc_state_field_type_31_is_repeated(
      control_io_metadata_init_bits_desc_state_field_type_31_is_repeated),
    .io_metadata_init_bits_desc_state_field_type_31_field_type(
      control_io_metadata_init_bits_desc_state_field_type_31_field_type),
    .io_metadata_init_bits_desc_state_field_type_31_sub_class_id(
      control_io_metadata_init_bits_desc_state_field_type_31_sub_class_id),
    .io_metadata_init_bits_desc_state_field_type_31_is_host(
      control_io_metadata_init_bits_desc_state_field_type_31_is_host),
    .io_metadata_init_bits_desc_state_field_type_32_is_repeated(
      control_io_metadata_init_bits_desc_state_field_type_32_is_repeated),
    .io_metadata_init_bits_desc_state_field_type_32_field_type(
      control_io_metadata_init_bits_desc_state_field_type_32_field_type),
    .io_metadata_init_bits_desc_state_field_type_32_sub_class_id(
      control_io_metadata_init_bits_desc_state_field_type_32_sub_class_id),
    .io_metadata_init_bits_desc_state_field_type_32_is_host(
      control_io_metadata_init_bits_desc_state_field_type_32_is_host),
    .io_ser_cmd_ready(control_io_ser_cmd_ready),
    .io_ser_cmd_valid(control_io_ser_cmd_valid),
    .io_ser_cmd_bits_class_id(control_io_ser_cmd_bits_class_id),
    .io_ser_cmd_bits_host_base_addr(control_io_ser_cmd_bits_host_base_addr)
  );
  ila_debug instIlaDbg ( // @[FpgaCloudSerHw.scala 166:40]
    .clk(instIlaDbg_clk),
    .data_1(instIlaDbg_data_1),
    .data_0(instIlaDbg_data_0)
  );
  assign io_cmacPin_tx_p = 4'h0;
  assign io_cmacPin_tx_n = 4'h0;
  assign io_cmacPin2_tx_p = 4'h0;
  assign io_cmacPin2_tx_n = 4'h0;
  assign io_ddrPort2_axi_aw_valid = 1'h0; // @[AXI.scala 198:49]
  assign io_ddrPort2_axi_aw_bits_addr = 34'h0; // @[Util.scala 13:40 Util.scala 13:40]
  assign io_ddrPort2_axi_aw_bits_burst = 2'h1; // @[AXI.scala 51:33]
  assign io_ddrPort2_axi_aw_bits_cache = 4'h0;
  assign io_ddrPort2_axi_aw_bits_id = 4'h0; // @[Util.scala 13:40 Util.scala 13:40]
  assign io_ddrPort2_axi_aw_bits_len = 8'h0; // @[Util.scala 13:40 Util.scala 13:40]
  assign io_ddrPort2_axi_aw_bits_lock = 1'h0;
  assign io_ddrPort2_axi_aw_bits_prot = 3'h0;
  assign io_ddrPort2_axi_aw_bits_qos = 4'h0;
  assign io_ddrPort2_axi_aw_bits_region = 4'h0;
  assign io_ddrPort2_axi_aw_bits_size = 3'h6; // @[AXI.scala 52:33]
  assign io_ddrPort2_axi_ar_valid = 1'h0; // @[AXI.scala 197:49]
  assign io_ddrPort2_axi_ar_bits_addr = 34'h0; // @[Util.scala 13:40 Util.scala 13:40]
  assign io_ddrPort2_axi_ar_bits_burst = 2'h1; // @[AXI.scala 51:33]
  assign io_ddrPort2_axi_ar_bits_cache = 4'h0;
  assign io_ddrPort2_axi_ar_bits_id = 4'h0; // @[Util.scala 13:40 Util.scala 13:40]
  assign io_ddrPort2_axi_ar_bits_len = 8'h0; // @[Util.scala 13:40 Util.scala 13:40]
  assign io_ddrPort2_axi_ar_bits_lock = 1'h0;
  assign io_ddrPort2_axi_ar_bits_prot = 3'h0;
  assign io_ddrPort2_axi_ar_bits_qos = 4'h0;
  assign io_ddrPort2_axi_ar_bits_region = 4'h0;
  assign io_ddrPort2_axi_ar_bits_size = 3'h6; // @[AXI.scala 52:33]
  assign io_ddrPort2_axi_w_valid = 1'h0; // @[AXI.scala 199:49]
  assign io_ddrPort2_axi_w_bits_data = 512'h0; // @[Util.scala 13:40 Util.scala 13:40]
  assign io_ddrPort2_axi_w_bits_last = 1'h0; // @[Util.scala 13:40 Util.scala 13:40]
  assign io_ddrPort2_axi_w_bits_strb = 64'hffffffffffffffff; // @[Util.scala 34:55]
  assign io_ddrPort2_axi_r_ready = 1'h0; // @[AXI.scala 200:49]
  assign io_ddrPort2_axi_b_ready = 1'h1; // @[AXI.scala 201:49]
  assign io_qdma_m_axib_awready = qdma_io_qdma_port_m_axib_awready; // @[FpgaCloudSerHw.scala 85:33]
  assign io_qdma_m_axib_wready = qdma_io_qdma_port_m_axib_wready; // @[FpgaCloudSerHw.scala 85:33]
  assign io_qdma_m_axib_bid = qdma_io_qdma_port_m_axib_bid; // @[FpgaCloudSerHw.scala 85:33]
  assign io_qdma_m_axib_bresp = qdma_io_qdma_port_m_axib_bresp; // @[FpgaCloudSerHw.scala 85:33]
  assign io_qdma_m_axib_bvalid = qdma_io_qdma_port_m_axib_bvalid; // @[FpgaCloudSerHw.scala 85:33]
  assign io_qdma_m_axib_arready = qdma_io_qdma_port_m_axib_arready; // @[FpgaCloudSerHw.scala 85:33]
  assign io_qdma_m_axib_rid = qdma_io_qdma_port_m_axib_rid; // @[FpgaCloudSerHw.scala 85:33]
  assign io_qdma_m_axib_rdata = qdma_io_qdma_port_m_axib_rdata; // @[FpgaCloudSerHw.scala 85:33]
  assign io_qdma_m_axib_rresp = qdma_io_qdma_port_m_axib_rresp; // @[FpgaCloudSerHw.scala 85:33]
  assign io_qdma_m_axib_rlast = qdma_io_qdma_port_m_axib_rlast; // @[FpgaCloudSerHw.scala 85:33]
  assign io_qdma_m_axib_rvalid = qdma_io_qdma_port_m_axib_rvalid; // @[FpgaCloudSerHw.scala 85:33]
  assign io_qdma_m_axil_awready = qdma_io_qdma_port_m_axil_awready; // @[FpgaCloudSerHw.scala 85:33]
  assign io_qdma_m_axil_wready = qdma_io_qdma_port_m_axil_wready; // @[FpgaCloudSerHw.scala 85:33]
  assign io_qdma_m_axil_bresp = qdma_io_qdma_port_m_axil_bresp; // @[FpgaCloudSerHw.scala 85:33]
  assign io_qdma_m_axil_bvalid = qdma_io_qdma_port_m_axil_bvalid; // @[FpgaCloudSerHw.scala 85:33]
  assign io_qdma_m_axil_arready = qdma_io_qdma_port_m_axil_arready; // @[FpgaCloudSerHw.scala 85:33]
  assign io_qdma_m_axil_rdata = qdma_io_qdma_port_m_axil_rdata; // @[FpgaCloudSerHw.scala 85:33]
  assign io_qdma_m_axil_rresp = qdma_io_qdma_port_m_axil_rresp; // @[FpgaCloudSerHw.scala 85:33]
  assign io_qdma_m_axil_rvalid = qdma_io_qdma_port_m_axil_rvalid; // @[FpgaCloudSerHw.scala 85:33]
  assign io_qdma_soft_reset_n = 1'h1; // @[FpgaCloudSerHw.scala 85:33]
  assign io_qdma_h2c_byp_in_st_addr = qdma_io_qdma_port_h2c_byp_in_st_addr; // @[FpgaCloudSerHw.scala 85:33]
  assign io_qdma_h2c_byp_in_st_len = qdma_io_qdma_port_h2c_byp_in_st_len; // @[FpgaCloudSerHw.scala 85:33]
  assign io_qdma_h2c_byp_in_st_eop = qdma_io_qdma_port_h2c_byp_in_st_eop; // @[FpgaCloudSerHw.scala 85:33]
  assign io_qdma_h2c_byp_in_st_sop = qdma_io_qdma_port_h2c_byp_in_st_sop; // @[FpgaCloudSerHw.scala 85:33]
  assign io_qdma_h2c_byp_in_st_mrkr_req = qdma_io_qdma_port_h2c_byp_in_st_mrkr_req; // @[FpgaCloudSerHw.scala 85:33]
  assign io_qdma_h2c_byp_in_st_sdi = qdma_io_qdma_port_h2c_byp_in_st_sdi; // @[FpgaCloudSerHw.scala 85:33]
  assign io_qdma_h2c_byp_in_st_qid = qdma_io_qdma_port_h2c_byp_in_st_qid; // @[FpgaCloudSerHw.scala 85:33]
  assign io_qdma_h2c_byp_in_st_error = qdma_io_qdma_port_h2c_byp_in_st_error; // @[FpgaCloudSerHw.scala 85:33]
  assign io_qdma_h2c_byp_in_st_func = qdma_io_qdma_port_h2c_byp_in_st_func; // @[FpgaCloudSerHw.scala 85:33]
  assign io_qdma_h2c_byp_in_st_cidx = qdma_io_qdma_port_h2c_byp_in_st_cidx; // @[FpgaCloudSerHw.scala 85:33]
  assign io_qdma_h2c_byp_in_st_port_id = qdma_io_qdma_port_h2c_byp_in_st_port_id; // @[FpgaCloudSerHw.scala 85:33]
  assign io_qdma_h2c_byp_in_st_no_dma = qdma_io_qdma_port_h2c_byp_in_st_no_dma; // @[FpgaCloudSerHw.scala 85:33]
  assign io_qdma_h2c_byp_in_st_vld = qdma_io_qdma_port_h2c_byp_in_st_vld; // @[FpgaCloudSerHw.scala 85:33]
  assign io_qdma_c2h_byp_in_st_csh_addr = qdma_io_qdma_port_c2h_byp_in_st_csh_addr; // @[FpgaCloudSerHw.scala 85:33]
  assign io_qdma_c2h_byp_in_st_csh_qid = qdma_io_qdma_port_c2h_byp_in_st_csh_qid; // @[FpgaCloudSerHw.scala 85:33]
  assign io_qdma_c2h_byp_in_st_csh_error = qdma_io_qdma_port_c2h_byp_in_st_csh_error; // @[FpgaCloudSerHw.scala 85:33]
  assign io_qdma_c2h_byp_in_st_csh_func = qdma_io_qdma_port_c2h_byp_in_st_csh_func; // @[FpgaCloudSerHw.scala 85:33]
  assign io_qdma_c2h_byp_in_st_csh_port_id = qdma_io_qdma_port_c2h_byp_in_st_csh_port_id; // @[FpgaCloudSerHw.scala 85:33]
  assign io_qdma_c2h_byp_in_st_csh_pfch_tag = qdma_io_qdma_port_c2h_byp_in_st_csh_pfch_tag; // @[FpgaCloudSerHw.scala 85:33]
  assign io_qdma_c2h_byp_in_st_csh_vld = qdma_io_qdma_port_c2h_byp_in_st_csh_vld; // @[FpgaCloudSerHw.scala 85:33]
  assign io_qdma_s_axis_c2h_tdata = qdma_io_qdma_port_s_axis_c2h_tdata; // @[FpgaCloudSerHw.scala 85:33]
  assign io_qdma_s_axis_c2h_tcrc = qdma_io_qdma_port_s_axis_c2h_tcrc; // @[FpgaCloudSerHw.scala 85:33]
  assign io_qdma_s_axis_c2h_ctrl_marker = qdma_io_qdma_port_s_axis_c2h_ctrl_marker; // @[FpgaCloudSerHw.scala 85:33]
  assign io_qdma_s_axis_c2h_ctrl_ecc = qdma_io_qdma_port_s_axis_c2h_ctrl_ecc; // @[FpgaCloudSerHw.scala 85:33]
  assign io_qdma_s_axis_c2h_ctrl_len = qdma_io_qdma_port_s_axis_c2h_ctrl_len; // @[FpgaCloudSerHw.scala 85:33]
  assign io_qdma_s_axis_c2h_ctrl_port_id = qdma_io_qdma_port_s_axis_c2h_ctrl_port_id; // @[FpgaCloudSerHw.scala 85:33]
  assign io_qdma_s_axis_c2h_ctrl_qid = qdma_io_qdma_port_s_axis_c2h_ctrl_qid; // @[FpgaCloudSerHw.scala 85:33]
  assign io_qdma_s_axis_c2h_ctrl_has_cmpt = qdma_io_qdma_port_s_axis_c2h_ctrl_has_cmpt; // @[FpgaCloudSerHw.scala 85:33]
  assign io_qdma_s_axis_c2h_mty = qdma_io_qdma_port_s_axis_c2h_mty; // @[FpgaCloudSerHw.scala 85:33]
  assign io_qdma_s_axis_c2h_tlast = qdma_io_qdma_port_s_axis_c2h_tlast; // @[FpgaCloudSerHw.scala 85:33]
  assign io_qdma_s_axis_c2h_tvalid = qdma_io_qdma_port_s_axis_c2h_tvalid; // @[FpgaCloudSerHw.scala 85:33]
  assign io_qdma_m_axis_h2c_tready = qdma_io_qdma_port_m_axis_h2c_tready; // @[FpgaCloudSerHw.scala 85:33]
  assign io_qdma_s_axis_c2h_cmpt_tdata = 512'h0; // @[FpgaCloudSerHw.scala 85:33]
  assign io_qdma_s_axis_c2h_cmpt_size = 2'h0; // @[FpgaCloudSerHw.scala 85:33]
  assign io_qdma_s_axis_c2h_cmpt_dpar = 16'h0; // @[FpgaCloudSerHw.scala 85:33]
  assign io_qdma_s_axis_c2h_cmpt_tvalid = 1'h0; // @[FpgaCloudSerHw.scala 85:33]
  assign io_qdma_s_axis_c2h_cmpt_ctrl_qid = 11'h0; // @[FpgaCloudSerHw.scala 85:33]
  assign io_qdma_s_axis_c2h_cmpt_ctrl_cmpt_type = 2'h0; // @[FpgaCloudSerHw.scala 85:33]
  assign io_qdma_s_axis_c2h_cmpt_ctrl_wait_pld_pkt_id = 16'h0; // @[FpgaCloudSerHw.scala 85:33]
  assign io_qdma_s_axis_c2h_cmpt_ctrl_no_wrb_marker = 1'h0; // @[FpgaCloudSerHw.scala 85:33]
  assign io_qdma_s_axis_c2h_cmpt_ctrl_port_id = 3'h0; // @[FpgaCloudSerHw.scala 85:33]
  assign io_qdma_s_axis_c2h_cmpt_ctrl_marker = 1'h0; // @[FpgaCloudSerHw.scala 85:33]
  assign io_qdma_s_axis_c2h_cmpt_ctrl_user_trig = 1'h0; // @[FpgaCloudSerHw.scala 85:33]
  assign io_qdma_s_axis_c2h_cmpt_ctrl_col_idx = 3'h0; // @[FpgaCloudSerHw.scala 85:33]
  assign io_qdma_s_axis_c2h_cmpt_ctrl_err_idx = 3'h0; // @[FpgaCloudSerHw.scala 85:33]
  assign io_qdma_h2c_byp_out_rdy = 1'h1; // @[FpgaCloudSerHw.scala 85:33]
  assign io_qdma_c2h_byp_out_rdy = 1'h1; // @[FpgaCloudSerHw.scala 85:33]
  assign io_qdma_tm_dsc_sts_rdy = 1'h1; // @[FpgaCloudSerHw.scala 85:33]
  assign io_qdma_dsc_crdt_in_vld = 1'h0; // @[FpgaCloudSerHw.scala 85:33]
  assign io_qdma_dsc_crdt_in_dir = 1'h0; // @[FpgaCloudSerHw.scala 85:33]
  assign io_qdma_dsc_crdt_in_fence = 1'h0; // @[FpgaCloudSerHw.scala 85:33]
  assign io_qdma_dsc_crdt_in_qid = 11'h0; // @[FpgaCloudSerHw.scala 85:33]
  assign io_qdma_dsc_crdt_in_crdt = 16'h0; // @[FpgaCloudSerHw.scala 85:33]
  assign io_qdma_qsts_out_rdy = 1'h1; // @[FpgaCloudSerHw.scala 85:33]
  assign io_qdma_usr_irq_in_vld = 1'h0; // @[FpgaCloudSerHw.scala 85:33]
  assign io_qdma_usr_irq_in_vec = 11'h0; // @[FpgaCloudSerHw.scala 85:33]
  assign io_qdma_usr_irq_in_fnc = 8'h0; // @[FpgaCloudSerHw.scala 85:33]
  assign S_BSCAN_tdo = dbgBridgeInst_S_BSCAN_tdo; // @[DebugBridge.scala 65:53]
  assign dbgBridgeInst_clk = clock; // @[DebugBridge.scala 59:49]
  assign dbgBridgeInst_S_BSCAN_drck = S_BSCAN_drck; // @[DebugBridge.scala 60:53]
  assign dbgBridgeInst_S_BSCAN_shift = S_BSCAN_shift; // @[DebugBridge.scala 61:53]
  assign dbgBridgeInst_S_BSCAN_tdi = S_BSCAN_tdi; // @[DebugBridge.scala 62:53]
  assign dbgBridgeInst_S_BSCAN_update = S_BSCAN_update; // @[DebugBridge.scala 63:53]
  assign dbgBridgeInst_S_BSCAN_sel = S_BSCAN_sel; // @[DebugBridge.scala 64:53]
  assign dbgBridgeInst_S_BSCAN_tms = S_BSCAN_tms; // @[DebugBridge.scala 66:53]
  assign dbgBridgeInst_S_BSCAN_tck = S_BSCAN_tck; // @[DebugBridge.scala 67:53]
  assign dbgBridgeInst_S_BSCAN_runtest = S_BSCAN_runtest; // @[DebugBridge.scala 68:53]
  assign dbgBridgeInst_S_BSCAN_reset = S_BSCAN_reset; // @[DebugBridge.scala 69:53]
  assign dbgBridgeInst_S_BSCAN_capture = S_BSCAN_capture; // @[DebugBridge.scala 70:53]
  assign dbgBridgeInst_S_BSCAN_bscanid_en = S_BSCAN_bscanid_en; // @[DebugBridge.scala 71:49]
  assign hbmDriver_clock = io_sysClk;
  assign qdma_io_qdma_port_axi_aclk = io_qdma_axi_aclk; // @[FpgaCloudSerHw.scala 85:33]
  assign qdma_io_qdma_port_axi_aresetn = io_qdma_axi_aresetn; // @[FpgaCloudSerHw.scala 85:33]
  assign qdma_io_qdma_port_m_axib_awid = io_qdma_m_axib_awid; // @[FpgaCloudSerHw.scala 85:33]
  assign qdma_io_qdma_port_m_axib_awaddr = io_qdma_m_axib_awaddr; // @[FpgaCloudSerHw.scala 85:33]
  assign qdma_io_qdma_port_m_axib_awlen = io_qdma_m_axib_awlen; // @[FpgaCloudSerHw.scala 85:33]
  assign qdma_io_qdma_port_m_axib_awsize = io_qdma_m_axib_awsize; // @[FpgaCloudSerHw.scala 85:33]
  assign qdma_io_qdma_port_m_axib_awburst = io_qdma_m_axib_awburst; // @[FpgaCloudSerHw.scala 85:33]
  assign qdma_io_qdma_port_m_axib_awprot = io_qdma_m_axib_awprot; // @[FpgaCloudSerHw.scala 85:33]
  assign qdma_io_qdma_port_m_axib_awlock = io_qdma_m_axib_awlock; // @[FpgaCloudSerHw.scala 85:33]
  assign qdma_io_qdma_port_m_axib_awcache = io_qdma_m_axib_awcache; // @[FpgaCloudSerHw.scala 85:33]
  assign qdma_io_qdma_port_m_axib_awvalid = io_qdma_m_axib_awvalid; // @[FpgaCloudSerHw.scala 85:33]
  assign qdma_io_qdma_port_m_axib_wdata = io_qdma_m_axib_wdata; // @[FpgaCloudSerHw.scala 85:33]
  assign qdma_io_qdma_port_m_axib_wstrb = io_qdma_m_axib_wstrb; // @[FpgaCloudSerHw.scala 85:33]
  assign qdma_io_qdma_port_m_axib_wlast = io_qdma_m_axib_wlast; // @[FpgaCloudSerHw.scala 85:33]
  assign qdma_io_qdma_port_m_axib_wvalid = io_qdma_m_axib_wvalid; // @[FpgaCloudSerHw.scala 85:33]
  assign qdma_io_qdma_port_m_axib_bready = io_qdma_m_axib_bready; // @[FpgaCloudSerHw.scala 85:33]
  assign qdma_io_qdma_port_m_axib_arid = io_qdma_m_axib_arid; // @[FpgaCloudSerHw.scala 85:33]
  assign qdma_io_qdma_port_m_axib_araddr = io_qdma_m_axib_araddr; // @[FpgaCloudSerHw.scala 85:33]
  assign qdma_io_qdma_port_m_axib_arlen = io_qdma_m_axib_arlen; // @[FpgaCloudSerHw.scala 85:33]
  assign qdma_io_qdma_port_m_axib_arsize = io_qdma_m_axib_arsize; // @[FpgaCloudSerHw.scala 85:33]
  assign qdma_io_qdma_port_m_axib_arburst = io_qdma_m_axib_arburst; // @[FpgaCloudSerHw.scala 85:33]
  assign qdma_io_qdma_port_m_axib_arprot = io_qdma_m_axib_arprot; // @[FpgaCloudSerHw.scala 85:33]
  assign qdma_io_qdma_port_m_axib_arlock = io_qdma_m_axib_arlock; // @[FpgaCloudSerHw.scala 85:33]
  assign qdma_io_qdma_port_m_axib_arcache = io_qdma_m_axib_arcache; // @[FpgaCloudSerHw.scala 85:33]
  assign qdma_io_qdma_port_m_axib_arvalid = io_qdma_m_axib_arvalid; // @[FpgaCloudSerHw.scala 85:33]
  assign qdma_io_qdma_port_m_axib_rready = io_qdma_m_axib_rready; // @[FpgaCloudSerHw.scala 85:33]
  assign qdma_io_qdma_port_m_axil_awaddr = io_qdma_m_axil_awaddr; // @[FpgaCloudSerHw.scala 85:33]
  assign qdma_io_qdma_port_m_axil_awvalid = io_qdma_m_axil_awvalid; // @[FpgaCloudSerHw.scala 85:33]
  assign qdma_io_qdma_port_m_axil_wdata = io_qdma_m_axil_wdata; // @[FpgaCloudSerHw.scala 85:33]
  assign qdma_io_qdma_port_m_axil_wstrb = io_qdma_m_axil_wstrb; // @[FpgaCloudSerHw.scala 85:33]
  assign qdma_io_qdma_port_m_axil_wvalid = io_qdma_m_axil_wvalid; // @[FpgaCloudSerHw.scala 85:33]
  assign qdma_io_qdma_port_m_axil_bready = io_qdma_m_axil_bready; // @[FpgaCloudSerHw.scala 85:33]
  assign qdma_io_qdma_port_m_axil_araddr = io_qdma_m_axil_araddr; // @[FpgaCloudSerHw.scala 85:33]
  assign qdma_io_qdma_port_m_axil_arvalid = io_qdma_m_axil_arvalid; // @[FpgaCloudSerHw.scala 85:33]
  assign qdma_io_qdma_port_m_axil_rready = io_qdma_m_axil_rready; // @[FpgaCloudSerHw.scala 85:33]
  assign qdma_io_qdma_port_h2c_byp_in_st_rdy = io_qdma_h2c_byp_in_st_rdy; // @[FpgaCloudSerHw.scala 85:33]
  assign qdma_io_qdma_port_c2h_byp_in_st_csh_rdy = io_qdma_c2h_byp_in_st_csh_rdy; // @[FpgaCloudSerHw.scala 85:33]
  assign qdma_io_qdma_port_s_axis_c2h_tready = io_qdma_s_axis_c2h_tready; // @[FpgaCloudSerHw.scala 85:33]
  assign qdma_io_qdma_port_m_axis_h2c_tdata = io_qdma_m_axis_h2c_tdata; // @[FpgaCloudSerHw.scala 85:33]
  assign qdma_io_qdma_port_m_axis_h2c_tcrc = io_qdma_m_axis_h2c_tcrc; // @[FpgaCloudSerHw.scala 85:33]
  assign qdma_io_qdma_port_m_axis_h2c_tuser_qid = io_qdma_m_axis_h2c_tuser_qid; // @[FpgaCloudSerHw.scala 85:33]
  assign qdma_io_qdma_port_m_axis_h2c_tuser_port_id = io_qdma_m_axis_h2c_tuser_port_id; // @[FpgaCloudSerHw.scala 85:33]
  assign qdma_io_qdma_port_m_axis_h2c_tuser_err = io_qdma_m_axis_h2c_tuser_err; // @[FpgaCloudSerHw.scala 85:33]
  assign qdma_io_qdma_port_m_axis_h2c_tuser_mdata = io_qdma_m_axis_h2c_tuser_mdata; // @[FpgaCloudSerHw.scala 85:33]
  assign qdma_io_qdma_port_m_axis_h2c_tuser_mty = io_qdma_m_axis_h2c_tuser_mty; // @[FpgaCloudSerHw.scala 85:33]
  assign qdma_io_qdma_port_m_axis_h2c_tuser_zero_byte = io_qdma_m_axis_h2c_tuser_zero_byte; // @[FpgaCloudSerHw.scala 85:33]
  assign qdma_io_qdma_port_m_axis_h2c_tlast = io_qdma_m_axis_h2c_tlast; // @[FpgaCloudSerHw.scala 85:33]
  assign qdma_io_qdma_port_m_axis_h2c_tvalid = io_qdma_m_axis_h2c_tvalid; // @[FpgaCloudSerHw.scala 85:33]
  assign qdma_io_user_clk = clock; // @[FpgaCloudSerHw.scala 61:31 FpgaCloudSerHw.scala 82:25]
  assign qdma_io_user_arstn = ~reset; // @[FpgaCloudSerHw.scala 87:36]
  assign qdma_io_h2c_cmd_valid = ser_io_host_data_cmd_valid; // @[FpgaCloudSerHw.scala 129:53]
  assign qdma_io_h2c_cmd_bits_addr = ser_io_host_data_cmd_bits_vaddr; // @[FpgaCloudSerHw.scala 131:53]
  assign qdma_io_h2c_cmd_bits_len = ser_io_host_data_cmd_bits_length; // @[FpgaCloudSerHw.scala 132:61]
  assign qdma_io_reg_status_300 = {{31'd0}, done_en}; // @[FpgaCloudSerHw.scala 180:49]
  assign qdma_io_reg_status_400 = qdma_io_tlb_miss_count; // @[Collector.scala 211:35]
  assign qdma_io_reg_status_401 = qdma_counter_0; // @[Collector.scala 211:35]
  assign qdma_io_reg_status_402 = qdma_counter_1_0; // @[Collector.scala 211:35]
  assign qdma_io_reg_status_403 = qdma_counter_2_1; // @[Collector.scala 211:35]
  assign qdma_io_reg_status_404 = qdma_counter_3_1; // @[Collector.scala 211:35]
  assign qdma_io_reg_status_405 = qdma_counter_4_0; // @[Collector.scala 211:35]
  assign qdma_io_reg_status_406 = qdma_counter_5_0; // @[Collector.scala 211:35]
  assign qdma_io_reg_status_407 = qdma_counter_6_0; // @[Collector.scala 211:35]
  assign qdma_io_reg_status_408 = qdma_counter_7_0; // @[Collector.scala 211:35]
  assign qdma_io_reg_status_409 = ser_counter_8; // @[Collector.scala 211:35]
  assign qdma_io_reg_status_410 = ser_counter_1_1; // @[Collector.scala 211:35]
  assign qdma_io_reg_status_411 = ser_counter_2_0; // @[Collector.scala 211:35]
  assign qdma_io_reg_status_412 = ser_counter_3_0; // @[Collector.scala 211:35]
  assign qdma_io_reg_status_413 = meta_table_counter_5; // @[Collector.scala 211:35]
  assign qdma_io_reg_status_414 = {16'h0,qdma_io_reg_status_414_lo}; // @[Collector.scala 237:73]
  assign qdma_io_axib_aw_ready = control_io_axi_aw_ready; // @[FpgaCloudSerHw.scala 112:57]
  assign qdma_io_axib_w_ready = control_io_axi_w_ready; // @[FpgaCloudSerHw.scala 112:57]
  assign qdma_io_axib_r_bits_data = control_io_axi_r_bits_data; // @[FpgaCloudSerHw.scala 112:57]
  assign ser_clock = clock;
  assign ser_reset = ~userRstn; // @[FpgaCloudSerHw.scala 101:33]
  assign ser_io_meta_in_valid = control_io_ser_cmd_valid; // @[FpgaCloudSerHw.scala 115:49]
  assign ser_io_meta_in_bits_class_id = control_io_ser_cmd_bits_class_id; // @[FpgaCloudSerHw.scala 115:49]
  assign ser_io_meta_in_bits_host_base_addr = control_io_ser_cmd_bits_host_base_addr; // @[FpgaCloudSerHw.scala 115:49]
  assign ser_io_host_data_in_valid = qdma_io_h2c_data_valid; // @[FpgaCloudSerHw.scala 139:53]
  assign ser_io_host_data_cmd_ready = qdma_io_h2c_cmd_ready; // @[FpgaCloudSerHw.scala 130:53]
  assign ser_io_class_meta_req_ready = meta_table_io_s_class_meta_req_ready; // @[FpgaCloudSerHw.scala 121:31]
  assign ser_io_class_meta_rsp_valid = meta_table_io_s_class_meta_rsp_valid; // @[FpgaCloudSerHw.scala 122:31]
  assign ser_io_class_meta_rsp_bits_class_meta_max_field_num =
    meta_table_io_s_class_meta_rsp_bits_class_meta_max_field_num; // @[FpgaCloudSerHw.scala 122:31]
  assign ser_io_class_meta_rsp_bits_class_meta_field_type_0_is_repeated =
    meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_0_is_repeated; // @[FpgaCloudSerHw.scala 122:31]
  assign ser_io_class_meta_rsp_bits_class_meta_field_type_0_field_type =
    meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_0_field_type; // @[FpgaCloudSerHw.scala 122:31]
  assign ser_io_class_meta_rsp_bits_class_meta_field_type_0_sub_class_id =
    meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_0_sub_class_id; // @[FpgaCloudSerHw.scala 122:31]
  assign ser_io_class_meta_rsp_bits_class_meta_field_type_1_is_repeated =
    meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_1_is_repeated; // @[FpgaCloudSerHw.scala 122:31]
  assign ser_io_class_meta_rsp_bits_class_meta_field_type_1_field_type =
    meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_1_field_type; // @[FpgaCloudSerHw.scala 122:31]
  assign ser_io_class_meta_rsp_bits_class_meta_field_type_1_sub_class_id =
    meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_1_sub_class_id; // @[FpgaCloudSerHw.scala 122:31]
  assign ser_io_class_meta_rsp_bits_class_meta_field_type_2_is_repeated =
    meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_2_is_repeated; // @[FpgaCloudSerHw.scala 122:31]
  assign ser_io_class_meta_rsp_bits_class_meta_field_type_2_field_type =
    meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_2_field_type; // @[FpgaCloudSerHw.scala 122:31]
  assign ser_io_class_meta_rsp_bits_class_meta_field_type_2_sub_class_id =
    meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_2_sub_class_id; // @[FpgaCloudSerHw.scala 122:31]
  assign ser_io_class_meta_rsp_bits_class_meta_field_type_3_is_repeated =
    meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_3_is_repeated; // @[FpgaCloudSerHw.scala 122:31]
  assign ser_io_class_meta_rsp_bits_class_meta_field_type_3_field_type =
    meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_3_field_type; // @[FpgaCloudSerHw.scala 122:31]
  assign ser_io_class_meta_rsp_bits_class_meta_field_type_3_sub_class_id =
    meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_3_sub_class_id; // @[FpgaCloudSerHw.scala 122:31]
  assign ser_io_class_meta_rsp_bits_class_meta_field_type_4_is_repeated =
    meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_4_is_repeated; // @[FpgaCloudSerHw.scala 122:31]
  assign ser_io_class_meta_rsp_bits_class_meta_field_type_4_field_type =
    meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_4_field_type; // @[FpgaCloudSerHw.scala 122:31]
  assign ser_io_class_meta_rsp_bits_class_meta_field_type_4_sub_class_id =
    meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_4_sub_class_id; // @[FpgaCloudSerHw.scala 122:31]
  assign ser_io_class_meta_rsp_bits_class_meta_field_type_5_is_repeated =
    meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_5_is_repeated; // @[FpgaCloudSerHw.scala 122:31]
  assign ser_io_class_meta_rsp_bits_class_meta_field_type_5_field_type =
    meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_5_field_type; // @[FpgaCloudSerHw.scala 122:31]
  assign ser_io_class_meta_rsp_bits_class_meta_field_type_5_sub_class_id =
    meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_5_sub_class_id; // @[FpgaCloudSerHw.scala 122:31]
  assign ser_io_class_meta_rsp_bits_class_meta_field_type_6_is_repeated =
    meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_6_is_repeated; // @[FpgaCloudSerHw.scala 122:31]
  assign ser_io_class_meta_rsp_bits_class_meta_field_type_6_field_type =
    meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_6_field_type; // @[FpgaCloudSerHw.scala 122:31]
  assign ser_io_class_meta_rsp_bits_class_meta_field_type_6_sub_class_id =
    meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_6_sub_class_id; // @[FpgaCloudSerHw.scala 122:31]
  assign ser_io_class_meta_rsp_bits_class_meta_field_type_7_is_repeated =
    meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_7_is_repeated; // @[FpgaCloudSerHw.scala 122:31]
  assign ser_io_class_meta_rsp_bits_class_meta_field_type_7_field_type =
    meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_7_field_type; // @[FpgaCloudSerHw.scala 122:31]
  assign ser_io_class_meta_rsp_bits_class_meta_field_type_7_sub_class_id =
    meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_7_sub_class_id; // @[FpgaCloudSerHw.scala 122:31]
  assign ser_io_class_meta_rsp_bits_class_meta_field_type_8_is_repeated =
    meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_8_is_repeated; // @[FpgaCloudSerHw.scala 122:31]
  assign ser_io_class_meta_rsp_bits_class_meta_field_type_8_field_type =
    meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_8_field_type; // @[FpgaCloudSerHw.scala 122:31]
  assign ser_io_class_meta_rsp_bits_class_meta_field_type_8_sub_class_id =
    meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_8_sub_class_id; // @[FpgaCloudSerHw.scala 122:31]
  assign ser_io_class_meta_rsp_bits_class_meta_field_type_9_is_repeated =
    meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_9_is_repeated; // @[FpgaCloudSerHw.scala 122:31]
  assign ser_io_class_meta_rsp_bits_class_meta_field_type_9_field_type =
    meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_9_field_type; // @[FpgaCloudSerHw.scala 122:31]
  assign ser_io_class_meta_rsp_bits_class_meta_field_type_9_sub_class_id =
    meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_9_sub_class_id; // @[FpgaCloudSerHw.scala 122:31]
  assign ser_io_class_meta_rsp_bits_class_meta_field_type_10_is_repeated =
    meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_10_is_repeated; // @[FpgaCloudSerHw.scala 122:31]
  assign ser_io_class_meta_rsp_bits_class_meta_field_type_10_field_type =
    meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_10_field_type; // @[FpgaCloudSerHw.scala 122:31]
  assign ser_io_class_meta_rsp_bits_class_meta_field_type_10_sub_class_id =
    meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_10_sub_class_id; // @[FpgaCloudSerHw.scala 122:31]
  assign ser_io_class_meta_rsp_bits_class_meta_field_type_11_is_repeated =
    meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_11_is_repeated; // @[FpgaCloudSerHw.scala 122:31]
  assign ser_io_class_meta_rsp_bits_class_meta_field_type_11_field_type =
    meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_11_field_type; // @[FpgaCloudSerHw.scala 122:31]
  assign ser_io_class_meta_rsp_bits_class_meta_field_type_11_sub_class_id =
    meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_11_sub_class_id; // @[FpgaCloudSerHw.scala 122:31]
  assign ser_io_class_meta_rsp_bits_class_meta_field_type_12_is_repeated =
    meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_12_is_repeated; // @[FpgaCloudSerHw.scala 122:31]
  assign ser_io_class_meta_rsp_bits_class_meta_field_type_12_field_type =
    meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_12_field_type; // @[FpgaCloudSerHw.scala 122:31]
  assign ser_io_class_meta_rsp_bits_class_meta_field_type_12_sub_class_id =
    meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_12_sub_class_id; // @[FpgaCloudSerHw.scala 122:31]
  assign ser_io_class_meta_rsp_bits_class_meta_field_type_13_is_repeated =
    meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_13_is_repeated; // @[FpgaCloudSerHw.scala 122:31]
  assign ser_io_class_meta_rsp_bits_class_meta_field_type_13_field_type =
    meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_13_field_type; // @[FpgaCloudSerHw.scala 122:31]
  assign ser_io_class_meta_rsp_bits_class_meta_field_type_13_sub_class_id =
    meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_13_sub_class_id; // @[FpgaCloudSerHw.scala 122:31]
  assign ser_io_class_meta_rsp_bits_class_meta_field_type_14_is_repeated =
    meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_14_is_repeated; // @[FpgaCloudSerHw.scala 122:31]
  assign ser_io_class_meta_rsp_bits_class_meta_field_type_14_field_type =
    meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_14_field_type; // @[FpgaCloudSerHw.scala 122:31]
  assign ser_io_class_meta_rsp_bits_class_meta_field_type_14_sub_class_id =
    meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_14_sub_class_id; // @[FpgaCloudSerHw.scala 122:31]
  assign ser_io_class_meta_rsp_bits_class_meta_field_type_15_is_repeated =
    meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_15_is_repeated; // @[FpgaCloudSerHw.scala 122:31]
  assign ser_io_class_meta_rsp_bits_class_meta_field_type_15_field_type =
    meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_15_field_type; // @[FpgaCloudSerHw.scala 122:31]
  assign ser_io_class_meta_rsp_bits_class_meta_field_type_15_sub_class_id =
    meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_15_sub_class_id; // @[FpgaCloudSerHw.scala 122:31]
  assign ser_io_class_meta_rsp_bits_class_meta_field_type_16_is_repeated =
    meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_16_is_repeated; // @[FpgaCloudSerHw.scala 122:31]
  assign ser_io_class_meta_rsp_bits_class_meta_field_type_16_field_type =
    meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_16_field_type; // @[FpgaCloudSerHw.scala 122:31]
  assign ser_io_class_meta_rsp_bits_class_meta_field_type_16_sub_class_id =
    meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_16_sub_class_id; // @[FpgaCloudSerHw.scala 122:31]
  assign ser_io_class_meta_rsp_bits_class_meta_field_type_17_is_repeated =
    meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_17_is_repeated; // @[FpgaCloudSerHw.scala 122:31]
  assign ser_io_class_meta_rsp_bits_class_meta_field_type_17_field_type =
    meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_17_field_type; // @[FpgaCloudSerHw.scala 122:31]
  assign ser_io_class_meta_rsp_bits_class_meta_field_type_17_sub_class_id =
    meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_17_sub_class_id; // @[FpgaCloudSerHw.scala 122:31]
  assign ser_io_class_meta_rsp_bits_class_meta_field_type_18_is_repeated =
    meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_18_is_repeated; // @[FpgaCloudSerHw.scala 122:31]
  assign ser_io_class_meta_rsp_bits_class_meta_field_type_18_field_type =
    meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_18_field_type; // @[FpgaCloudSerHw.scala 122:31]
  assign ser_io_class_meta_rsp_bits_class_meta_field_type_18_sub_class_id =
    meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_18_sub_class_id; // @[FpgaCloudSerHw.scala 122:31]
  assign ser_io_class_meta_rsp_bits_class_meta_field_type_19_is_repeated =
    meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_19_is_repeated; // @[FpgaCloudSerHw.scala 122:31]
  assign ser_io_class_meta_rsp_bits_class_meta_field_type_19_field_type =
    meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_19_field_type; // @[FpgaCloudSerHw.scala 122:31]
  assign ser_io_class_meta_rsp_bits_class_meta_field_type_19_sub_class_id =
    meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_19_sub_class_id; // @[FpgaCloudSerHw.scala 122:31]
  assign ser_io_class_meta_rsp_bits_class_meta_field_type_20_is_repeated =
    meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_20_is_repeated; // @[FpgaCloudSerHw.scala 122:31]
  assign ser_io_class_meta_rsp_bits_class_meta_field_type_20_field_type =
    meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_20_field_type; // @[FpgaCloudSerHw.scala 122:31]
  assign ser_io_class_meta_rsp_bits_class_meta_field_type_20_sub_class_id =
    meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_20_sub_class_id; // @[FpgaCloudSerHw.scala 122:31]
  assign ser_io_class_meta_rsp_bits_class_meta_field_type_21_is_repeated =
    meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_21_is_repeated; // @[FpgaCloudSerHw.scala 122:31]
  assign ser_io_class_meta_rsp_bits_class_meta_field_type_21_field_type =
    meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_21_field_type; // @[FpgaCloudSerHw.scala 122:31]
  assign ser_io_class_meta_rsp_bits_class_meta_field_type_21_sub_class_id =
    meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_21_sub_class_id; // @[FpgaCloudSerHw.scala 122:31]
  assign ser_io_class_meta_rsp_bits_class_meta_field_type_22_is_repeated =
    meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_22_is_repeated; // @[FpgaCloudSerHw.scala 122:31]
  assign ser_io_class_meta_rsp_bits_class_meta_field_type_22_field_type =
    meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_22_field_type; // @[FpgaCloudSerHw.scala 122:31]
  assign ser_io_class_meta_rsp_bits_class_meta_field_type_22_sub_class_id =
    meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_22_sub_class_id; // @[FpgaCloudSerHw.scala 122:31]
  assign ser_io_class_meta_rsp_bits_class_meta_field_type_23_is_repeated =
    meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_23_is_repeated; // @[FpgaCloudSerHw.scala 122:31]
  assign ser_io_class_meta_rsp_bits_class_meta_field_type_23_field_type =
    meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_23_field_type; // @[FpgaCloudSerHw.scala 122:31]
  assign ser_io_class_meta_rsp_bits_class_meta_field_type_23_sub_class_id =
    meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_23_sub_class_id; // @[FpgaCloudSerHw.scala 122:31]
  assign ser_io_class_meta_rsp_bits_class_meta_field_type_24_is_repeated =
    meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_24_is_repeated; // @[FpgaCloudSerHw.scala 122:31]
  assign ser_io_class_meta_rsp_bits_class_meta_field_type_24_field_type =
    meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_24_field_type; // @[FpgaCloudSerHw.scala 122:31]
  assign ser_io_class_meta_rsp_bits_class_meta_field_type_24_sub_class_id =
    meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_24_sub_class_id; // @[FpgaCloudSerHw.scala 122:31]
  assign ser_io_class_meta_rsp_bits_class_meta_field_type_25_is_repeated =
    meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_25_is_repeated; // @[FpgaCloudSerHw.scala 122:31]
  assign ser_io_class_meta_rsp_bits_class_meta_field_type_25_field_type =
    meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_25_field_type; // @[FpgaCloudSerHw.scala 122:31]
  assign ser_io_class_meta_rsp_bits_class_meta_field_type_25_sub_class_id =
    meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_25_sub_class_id; // @[FpgaCloudSerHw.scala 122:31]
  assign ser_io_class_meta_rsp_bits_class_meta_field_type_26_is_repeated =
    meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_26_is_repeated; // @[FpgaCloudSerHw.scala 122:31]
  assign ser_io_class_meta_rsp_bits_class_meta_field_type_26_field_type =
    meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_26_field_type; // @[FpgaCloudSerHw.scala 122:31]
  assign ser_io_class_meta_rsp_bits_class_meta_field_type_26_sub_class_id =
    meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_26_sub_class_id; // @[FpgaCloudSerHw.scala 122:31]
  assign ser_io_class_meta_rsp_bits_class_meta_field_type_27_is_repeated =
    meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_27_is_repeated; // @[FpgaCloudSerHw.scala 122:31]
  assign ser_io_class_meta_rsp_bits_class_meta_field_type_27_field_type =
    meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_27_field_type; // @[FpgaCloudSerHw.scala 122:31]
  assign ser_io_class_meta_rsp_bits_class_meta_field_type_27_sub_class_id =
    meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_27_sub_class_id; // @[FpgaCloudSerHw.scala 122:31]
  assign ser_io_class_meta_rsp_bits_class_meta_field_type_28_is_repeated =
    meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_28_is_repeated; // @[FpgaCloudSerHw.scala 122:31]
  assign ser_io_class_meta_rsp_bits_class_meta_field_type_28_field_type =
    meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_28_field_type; // @[FpgaCloudSerHw.scala 122:31]
  assign ser_io_class_meta_rsp_bits_class_meta_field_type_28_sub_class_id =
    meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_28_sub_class_id; // @[FpgaCloudSerHw.scala 122:31]
  assign ser_io_class_meta_rsp_bits_class_meta_field_type_29_is_repeated =
    meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_29_is_repeated; // @[FpgaCloudSerHw.scala 122:31]
  assign ser_io_class_meta_rsp_bits_class_meta_field_type_29_field_type =
    meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_29_field_type; // @[FpgaCloudSerHw.scala 122:31]
  assign ser_io_class_meta_rsp_bits_class_meta_field_type_29_sub_class_id =
    meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_29_sub_class_id; // @[FpgaCloudSerHw.scala 122:31]
  assign ser_io_class_meta_rsp_bits_class_meta_field_type_30_is_repeated =
    meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_30_is_repeated; // @[FpgaCloudSerHw.scala 122:31]
  assign ser_io_class_meta_rsp_bits_class_meta_field_type_30_field_type =
    meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_30_field_type; // @[FpgaCloudSerHw.scala 122:31]
  assign ser_io_class_meta_rsp_bits_class_meta_field_type_30_sub_class_id =
    meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_30_sub_class_id; // @[FpgaCloudSerHw.scala 122:31]
  assign ser_io_class_meta_rsp_bits_class_meta_field_type_31_is_repeated =
    meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_31_is_repeated; // @[FpgaCloudSerHw.scala 122:31]
  assign ser_io_class_meta_rsp_bits_class_meta_field_type_31_field_type =
    meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_31_field_type; // @[FpgaCloudSerHw.scala 122:31]
  assign ser_io_class_meta_rsp_bits_class_meta_field_type_31_sub_class_id =
    meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_31_sub_class_id; // @[FpgaCloudSerHw.scala 122:31]
  assign ser_io_class_meta_rsp_bits_class_meta_field_type_32_is_repeated =
    meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_32_is_repeated; // @[FpgaCloudSerHw.scala 122:31]
  assign ser_io_class_meta_rsp_bits_class_meta_field_type_32_field_type =
    meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_32_field_type; // @[FpgaCloudSerHw.scala 122:31]
  assign ser_io_class_meta_rsp_bits_class_meta_field_type_32_sub_class_id =
    meta_table_io_s_class_meta_rsp_bits_class_meta_field_type_32_sub_class_id; // @[FpgaCloudSerHw.scala 122:31]
  assign ser_io_done_ready = 1'h1; // @[FpgaCloudSerHw.scala 119:41]
  assign meta_table_clock = clock;
  assign meta_table_reset = ~userRstn; // @[FpgaCloudSerHw.scala 101:33]
  assign meta_table_io_class_meta_init_valid = control_io_metadata_init_valid; // @[FpgaCloudSerHw.scala 114:49]
  assign meta_table_io_class_meta_init_bits_class_id = control_io_metadata_init_bits_class_id; // @[FpgaCloudSerHw.scala 114:49]
  assign meta_table_io_class_meta_init_bits_desc_state_class_length =
    control_io_metadata_init_bits_desc_state_class_length; // @[FpgaCloudSerHw.scala 114:49]
  assign meta_table_io_class_meta_init_bits_desc_state_max_field_num =
    control_io_metadata_init_bits_desc_state_max_field_num; // @[FpgaCloudSerHw.scala 114:49]
  assign meta_table_io_class_meta_init_bits_desc_state_field_type_0_is_repeated =
    control_io_metadata_init_bits_desc_state_field_type_0_is_repeated; // @[FpgaCloudSerHw.scala 114:49]
  assign meta_table_io_class_meta_init_bits_desc_state_field_type_0_field_type =
    control_io_metadata_init_bits_desc_state_field_type_0_field_type; // @[FpgaCloudSerHw.scala 114:49]
  assign meta_table_io_class_meta_init_bits_desc_state_field_type_0_sub_class_id =
    control_io_metadata_init_bits_desc_state_field_type_0_sub_class_id; // @[FpgaCloudSerHw.scala 114:49]
  assign meta_table_io_class_meta_init_bits_desc_state_field_type_0_is_host =
    control_io_metadata_init_bits_desc_state_field_type_0_is_host; // @[FpgaCloudSerHw.scala 114:49]
  assign meta_table_io_class_meta_init_bits_desc_state_field_type_1_is_repeated =
    control_io_metadata_init_bits_desc_state_field_type_1_is_repeated; // @[FpgaCloudSerHw.scala 114:49]
  assign meta_table_io_class_meta_init_bits_desc_state_field_type_1_field_type =
    control_io_metadata_init_bits_desc_state_field_type_1_field_type; // @[FpgaCloudSerHw.scala 114:49]
  assign meta_table_io_class_meta_init_bits_desc_state_field_type_1_sub_class_id =
    control_io_metadata_init_bits_desc_state_field_type_1_sub_class_id; // @[FpgaCloudSerHw.scala 114:49]
  assign meta_table_io_class_meta_init_bits_desc_state_field_type_1_is_host =
    control_io_metadata_init_bits_desc_state_field_type_1_is_host; // @[FpgaCloudSerHw.scala 114:49]
  assign meta_table_io_class_meta_init_bits_desc_state_field_type_2_is_repeated =
    control_io_metadata_init_bits_desc_state_field_type_2_is_repeated; // @[FpgaCloudSerHw.scala 114:49]
  assign meta_table_io_class_meta_init_bits_desc_state_field_type_2_field_type =
    control_io_metadata_init_bits_desc_state_field_type_2_field_type; // @[FpgaCloudSerHw.scala 114:49]
  assign meta_table_io_class_meta_init_bits_desc_state_field_type_2_sub_class_id =
    control_io_metadata_init_bits_desc_state_field_type_2_sub_class_id; // @[FpgaCloudSerHw.scala 114:49]
  assign meta_table_io_class_meta_init_bits_desc_state_field_type_2_is_host =
    control_io_metadata_init_bits_desc_state_field_type_2_is_host; // @[FpgaCloudSerHw.scala 114:49]
  assign meta_table_io_class_meta_init_bits_desc_state_field_type_3_is_repeated =
    control_io_metadata_init_bits_desc_state_field_type_3_is_repeated; // @[FpgaCloudSerHw.scala 114:49]
  assign meta_table_io_class_meta_init_bits_desc_state_field_type_3_field_type =
    control_io_metadata_init_bits_desc_state_field_type_3_field_type; // @[FpgaCloudSerHw.scala 114:49]
  assign meta_table_io_class_meta_init_bits_desc_state_field_type_3_sub_class_id =
    control_io_metadata_init_bits_desc_state_field_type_3_sub_class_id; // @[FpgaCloudSerHw.scala 114:49]
  assign meta_table_io_class_meta_init_bits_desc_state_field_type_3_is_host =
    control_io_metadata_init_bits_desc_state_field_type_3_is_host; // @[FpgaCloudSerHw.scala 114:49]
  assign meta_table_io_class_meta_init_bits_desc_state_field_type_4_is_repeated =
    control_io_metadata_init_bits_desc_state_field_type_4_is_repeated; // @[FpgaCloudSerHw.scala 114:49]
  assign meta_table_io_class_meta_init_bits_desc_state_field_type_4_field_type =
    control_io_metadata_init_bits_desc_state_field_type_4_field_type; // @[FpgaCloudSerHw.scala 114:49]
  assign meta_table_io_class_meta_init_bits_desc_state_field_type_4_sub_class_id =
    control_io_metadata_init_bits_desc_state_field_type_4_sub_class_id; // @[FpgaCloudSerHw.scala 114:49]
  assign meta_table_io_class_meta_init_bits_desc_state_field_type_4_is_host =
    control_io_metadata_init_bits_desc_state_field_type_4_is_host; // @[FpgaCloudSerHw.scala 114:49]
  assign meta_table_io_class_meta_init_bits_desc_state_field_type_5_is_repeated =
    control_io_metadata_init_bits_desc_state_field_type_5_is_repeated; // @[FpgaCloudSerHw.scala 114:49]
  assign meta_table_io_class_meta_init_bits_desc_state_field_type_5_field_type =
    control_io_metadata_init_bits_desc_state_field_type_5_field_type; // @[FpgaCloudSerHw.scala 114:49]
  assign meta_table_io_class_meta_init_bits_desc_state_field_type_5_sub_class_id =
    control_io_metadata_init_bits_desc_state_field_type_5_sub_class_id; // @[FpgaCloudSerHw.scala 114:49]
  assign meta_table_io_class_meta_init_bits_desc_state_field_type_5_is_host =
    control_io_metadata_init_bits_desc_state_field_type_5_is_host; // @[FpgaCloudSerHw.scala 114:49]
  assign meta_table_io_class_meta_init_bits_desc_state_field_type_6_is_repeated =
    control_io_metadata_init_bits_desc_state_field_type_6_is_repeated; // @[FpgaCloudSerHw.scala 114:49]
  assign meta_table_io_class_meta_init_bits_desc_state_field_type_6_field_type =
    control_io_metadata_init_bits_desc_state_field_type_6_field_type; // @[FpgaCloudSerHw.scala 114:49]
  assign meta_table_io_class_meta_init_bits_desc_state_field_type_6_sub_class_id =
    control_io_metadata_init_bits_desc_state_field_type_6_sub_class_id; // @[FpgaCloudSerHw.scala 114:49]
  assign meta_table_io_class_meta_init_bits_desc_state_field_type_6_is_host =
    control_io_metadata_init_bits_desc_state_field_type_6_is_host; // @[FpgaCloudSerHw.scala 114:49]
  assign meta_table_io_class_meta_init_bits_desc_state_field_type_7_is_repeated =
    control_io_metadata_init_bits_desc_state_field_type_7_is_repeated; // @[FpgaCloudSerHw.scala 114:49]
  assign meta_table_io_class_meta_init_bits_desc_state_field_type_7_field_type =
    control_io_metadata_init_bits_desc_state_field_type_7_field_type; // @[FpgaCloudSerHw.scala 114:49]
  assign meta_table_io_class_meta_init_bits_desc_state_field_type_7_sub_class_id =
    control_io_metadata_init_bits_desc_state_field_type_7_sub_class_id; // @[FpgaCloudSerHw.scala 114:49]
  assign meta_table_io_class_meta_init_bits_desc_state_field_type_7_is_host =
    control_io_metadata_init_bits_desc_state_field_type_7_is_host; // @[FpgaCloudSerHw.scala 114:49]
  assign meta_table_io_class_meta_init_bits_desc_state_field_type_8_is_repeated =
    control_io_metadata_init_bits_desc_state_field_type_8_is_repeated; // @[FpgaCloudSerHw.scala 114:49]
  assign meta_table_io_class_meta_init_bits_desc_state_field_type_8_field_type =
    control_io_metadata_init_bits_desc_state_field_type_8_field_type; // @[FpgaCloudSerHw.scala 114:49]
  assign meta_table_io_class_meta_init_bits_desc_state_field_type_8_sub_class_id =
    control_io_metadata_init_bits_desc_state_field_type_8_sub_class_id; // @[FpgaCloudSerHw.scala 114:49]
  assign meta_table_io_class_meta_init_bits_desc_state_field_type_8_is_host =
    control_io_metadata_init_bits_desc_state_field_type_8_is_host; // @[FpgaCloudSerHw.scala 114:49]
  assign meta_table_io_class_meta_init_bits_desc_state_field_type_9_is_repeated =
    control_io_metadata_init_bits_desc_state_field_type_9_is_repeated; // @[FpgaCloudSerHw.scala 114:49]
  assign meta_table_io_class_meta_init_bits_desc_state_field_type_9_field_type =
    control_io_metadata_init_bits_desc_state_field_type_9_field_type; // @[FpgaCloudSerHw.scala 114:49]
  assign meta_table_io_class_meta_init_bits_desc_state_field_type_9_sub_class_id =
    control_io_metadata_init_bits_desc_state_field_type_9_sub_class_id; // @[FpgaCloudSerHw.scala 114:49]
  assign meta_table_io_class_meta_init_bits_desc_state_field_type_9_is_host =
    control_io_metadata_init_bits_desc_state_field_type_9_is_host; // @[FpgaCloudSerHw.scala 114:49]
  assign meta_table_io_class_meta_init_bits_desc_state_field_type_10_is_repeated =
    control_io_metadata_init_bits_desc_state_field_type_10_is_repeated; // @[FpgaCloudSerHw.scala 114:49]
  assign meta_table_io_class_meta_init_bits_desc_state_field_type_10_field_type =
    control_io_metadata_init_bits_desc_state_field_type_10_field_type; // @[FpgaCloudSerHw.scala 114:49]
  assign meta_table_io_class_meta_init_bits_desc_state_field_type_10_sub_class_id =
    control_io_metadata_init_bits_desc_state_field_type_10_sub_class_id; // @[FpgaCloudSerHw.scala 114:49]
  assign meta_table_io_class_meta_init_bits_desc_state_field_type_10_is_host =
    control_io_metadata_init_bits_desc_state_field_type_10_is_host; // @[FpgaCloudSerHw.scala 114:49]
  assign meta_table_io_class_meta_init_bits_desc_state_field_type_11_is_repeated =
    control_io_metadata_init_bits_desc_state_field_type_11_is_repeated; // @[FpgaCloudSerHw.scala 114:49]
  assign meta_table_io_class_meta_init_bits_desc_state_field_type_11_field_type =
    control_io_metadata_init_bits_desc_state_field_type_11_field_type; // @[FpgaCloudSerHw.scala 114:49]
  assign meta_table_io_class_meta_init_bits_desc_state_field_type_11_sub_class_id =
    control_io_metadata_init_bits_desc_state_field_type_11_sub_class_id; // @[FpgaCloudSerHw.scala 114:49]
  assign meta_table_io_class_meta_init_bits_desc_state_field_type_11_is_host =
    control_io_metadata_init_bits_desc_state_field_type_11_is_host; // @[FpgaCloudSerHw.scala 114:49]
  assign meta_table_io_class_meta_init_bits_desc_state_field_type_12_is_repeated =
    control_io_metadata_init_bits_desc_state_field_type_12_is_repeated; // @[FpgaCloudSerHw.scala 114:49]
  assign meta_table_io_class_meta_init_bits_desc_state_field_type_12_field_type =
    control_io_metadata_init_bits_desc_state_field_type_12_field_type; // @[FpgaCloudSerHw.scala 114:49]
  assign meta_table_io_class_meta_init_bits_desc_state_field_type_12_sub_class_id =
    control_io_metadata_init_bits_desc_state_field_type_12_sub_class_id; // @[FpgaCloudSerHw.scala 114:49]
  assign meta_table_io_class_meta_init_bits_desc_state_field_type_12_is_host =
    control_io_metadata_init_bits_desc_state_field_type_12_is_host; // @[FpgaCloudSerHw.scala 114:49]
  assign meta_table_io_class_meta_init_bits_desc_state_field_type_13_is_repeated =
    control_io_metadata_init_bits_desc_state_field_type_13_is_repeated; // @[FpgaCloudSerHw.scala 114:49]
  assign meta_table_io_class_meta_init_bits_desc_state_field_type_13_field_type =
    control_io_metadata_init_bits_desc_state_field_type_13_field_type; // @[FpgaCloudSerHw.scala 114:49]
  assign meta_table_io_class_meta_init_bits_desc_state_field_type_13_sub_class_id =
    control_io_metadata_init_bits_desc_state_field_type_13_sub_class_id; // @[FpgaCloudSerHw.scala 114:49]
  assign meta_table_io_class_meta_init_bits_desc_state_field_type_13_is_host =
    control_io_metadata_init_bits_desc_state_field_type_13_is_host; // @[FpgaCloudSerHw.scala 114:49]
  assign meta_table_io_class_meta_init_bits_desc_state_field_type_14_is_repeated =
    control_io_metadata_init_bits_desc_state_field_type_14_is_repeated; // @[FpgaCloudSerHw.scala 114:49]
  assign meta_table_io_class_meta_init_bits_desc_state_field_type_14_field_type =
    control_io_metadata_init_bits_desc_state_field_type_14_field_type; // @[FpgaCloudSerHw.scala 114:49]
  assign meta_table_io_class_meta_init_bits_desc_state_field_type_14_sub_class_id =
    control_io_metadata_init_bits_desc_state_field_type_14_sub_class_id; // @[FpgaCloudSerHw.scala 114:49]
  assign meta_table_io_class_meta_init_bits_desc_state_field_type_14_is_host =
    control_io_metadata_init_bits_desc_state_field_type_14_is_host; // @[FpgaCloudSerHw.scala 114:49]
  assign meta_table_io_class_meta_init_bits_desc_state_field_type_15_is_repeated =
    control_io_metadata_init_bits_desc_state_field_type_15_is_repeated; // @[FpgaCloudSerHw.scala 114:49]
  assign meta_table_io_class_meta_init_bits_desc_state_field_type_15_field_type =
    control_io_metadata_init_bits_desc_state_field_type_15_field_type; // @[FpgaCloudSerHw.scala 114:49]
  assign meta_table_io_class_meta_init_bits_desc_state_field_type_15_sub_class_id =
    control_io_metadata_init_bits_desc_state_field_type_15_sub_class_id; // @[FpgaCloudSerHw.scala 114:49]
  assign meta_table_io_class_meta_init_bits_desc_state_field_type_15_is_host =
    control_io_metadata_init_bits_desc_state_field_type_15_is_host; // @[FpgaCloudSerHw.scala 114:49]
  assign meta_table_io_class_meta_init_bits_desc_state_field_type_16_is_repeated =
    control_io_metadata_init_bits_desc_state_field_type_16_is_repeated; // @[FpgaCloudSerHw.scala 114:49]
  assign meta_table_io_class_meta_init_bits_desc_state_field_type_16_field_type =
    control_io_metadata_init_bits_desc_state_field_type_16_field_type; // @[FpgaCloudSerHw.scala 114:49]
  assign meta_table_io_class_meta_init_bits_desc_state_field_type_16_sub_class_id =
    control_io_metadata_init_bits_desc_state_field_type_16_sub_class_id; // @[FpgaCloudSerHw.scala 114:49]
  assign meta_table_io_class_meta_init_bits_desc_state_field_type_16_is_host =
    control_io_metadata_init_bits_desc_state_field_type_16_is_host; // @[FpgaCloudSerHw.scala 114:49]
  assign meta_table_io_class_meta_init_bits_desc_state_field_type_17_is_repeated =
    control_io_metadata_init_bits_desc_state_field_type_17_is_repeated; // @[FpgaCloudSerHw.scala 114:49]
  assign meta_table_io_class_meta_init_bits_desc_state_field_type_17_field_type =
    control_io_metadata_init_bits_desc_state_field_type_17_field_type; // @[FpgaCloudSerHw.scala 114:49]
  assign meta_table_io_class_meta_init_bits_desc_state_field_type_17_sub_class_id =
    control_io_metadata_init_bits_desc_state_field_type_17_sub_class_id; // @[FpgaCloudSerHw.scala 114:49]
  assign meta_table_io_class_meta_init_bits_desc_state_field_type_17_is_host =
    control_io_metadata_init_bits_desc_state_field_type_17_is_host; // @[FpgaCloudSerHw.scala 114:49]
  assign meta_table_io_class_meta_init_bits_desc_state_field_type_18_is_repeated =
    control_io_metadata_init_bits_desc_state_field_type_18_is_repeated; // @[FpgaCloudSerHw.scala 114:49]
  assign meta_table_io_class_meta_init_bits_desc_state_field_type_18_field_type =
    control_io_metadata_init_bits_desc_state_field_type_18_field_type; // @[FpgaCloudSerHw.scala 114:49]
  assign meta_table_io_class_meta_init_bits_desc_state_field_type_18_sub_class_id =
    control_io_metadata_init_bits_desc_state_field_type_18_sub_class_id; // @[FpgaCloudSerHw.scala 114:49]
  assign meta_table_io_class_meta_init_bits_desc_state_field_type_18_is_host =
    control_io_metadata_init_bits_desc_state_field_type_18_is_host; // @[FpgaCloudSerHw.scala 114:49]
  assign meta_table_io_class_meta_init_bits_desc_state_field_type_19_is_repeated =
    control_io_metadata_init_bits_desc_state_field_type_19_is_repeated; // @[FpgaCloudSerHw.scala 114:49]
  assign meta_table_io_class_meta_init_bits_desc_state_field_type_19_field_type =
    control_io_metadata_init_bits_desc_state_field_type_19_field_type; // @[FpgaCloudSerHw.scala 114:49]
  assign meta_table_io_class_meta_init_bits_desc_state_field_type_19_sub_class_id =
    control_io_metadata_init_bits_desc_state_field_type_19_sub_class_id; // @[FpgaCloudSerHw.scala 114:49]
  assign meta_table_io_class_meta_init_bits_desc_state_field_type_19_is_host =
    control_io_metadata_init_bits_desc_state_field_type_19_is_host; // @[FpgaCloudSerHw.scala 114:49]
  assign meta_table_io_class_meta_init_bits_desc_state_field_type_20_is_repeated =
    control_io_metadata_init_bits_desc_state_field_type_20_is_repeated; // @[FpgaCloudSerHw.scala 114:49]
  assign meta_table_io_class_meta_init_bits_desc_state_field_type_20_field_type =
    control_io_metadata_init_bits_desc_state_field_type_20_field_type; // @[FpgaCloudSerHw.scala 114:49]
  assign meta_table_io_class_meta_init_bits_desc_state_field_type_20_sub_class_id =
    control_io_metadata_init_bits_desc_state_field_type_20_sub_class_id; // @[FpgaCloudSerHw.scala 114:49]
  assign meta_table_io_class_meta_init_bits_desc_state_field_type_20_is_host =
    control_io_metadata_init_bits_desc_state_field_type_20_is_host; // @[FpgaCloudSerHw.scala 114:49]
  assign meta_table_io_class_meta_init_bits_desc_state_field_type_21_is_repeated =
    control_io_metadata_init_bits_desc_state_field_type_21_is_repeated; // @[FpgaCloudSerHw.scala 114:49]
  assign meta_table_io_class_meta_init_bits_desc_state_field_type_21_field_type =
    control_io_metadata_init_bits_desc_state_field_type_21_field_type; // @[FpgaCloudSerHw.scala 114:49]
  assign meta_table_io_class_meta_init_bits_desc_state_field_type_21_sub_class_id =
    control_io_metadata_init_bits_desc_state_field_type_21_sub_class_id; // @[FpgaCloudSerHw.scala 114:49]
  assign meta_table_io_class_meta_init_bits_desc_state_field_type_21_is_host =
    control_io_metadata_init_bits_desc_state_field_type_21_is_host; // @[FpgaCloudSerHw.scala 114:49]
  assign meta_table_io_class_meta_init_bits_desc_state_field_type_22_is_repeated =
    control_io_metadata_init_bits_desc_state_field_type_22_is_repeated; // @[FpgaCloudSerHw.scala 114:49]
  assign meta_table_io_class_meta_init_bits_desc_state_field_type_22_field_type =
    control_io_metadata_init_bits_desc_state_field_type_22_field_type; // @[FpgaCloudSerHw.scala 114:49]
  assign meta_table_io_class_meta_init_bits_desc_state_field_type_22_sub_class_id =
    control_io_metadata_init_bits_desc_state_field_type_22_sub_class_id; // @[FpgaCloudSerHw.scala 114:49]
  assign meta_table_io_class_meta_init_bits_desc_state_field_type_22_is_host =
    control_io_metadata_init_bits_desc_state_field_type_22_is_host; // @[FpgaCloudSerHw.scala 114:49]
  assign meta_table_io_class_meta_init_bits_desc_state_field_type_23_is_repeated =
    control_io_metadata_init_bits_desc_state_field_type_23_is_repeated; // @[FpgaCloudSerHw.scala 114:49]
  assign meta_table_io_class_meta_init_bits_desc_state_field_type_23_field_type =
    control_io_metadata_init_bits_desc_state_field_type_23_field_type; // @[FpgaCloudSerHw.scala 114:49]
  assign meta_table_io_class_meta_init_bits_desc_state_field_type_23_sub_class_id =
    control_io_metadata_init_bits_desc_state_field_type_23_sub_class_id; // @[FpgaCloudSerHw.scala 114:49]
  assign meta_table_io_class_meta_init_bits_desc_state_field_type_23_is_host =
    control_io_metadata_init_bits_desc_state_field_type_23_is_host; // @[FpgaCloudSerHw.scala 114:49]
  assign meta_table_io_class_meta_init_bits_desc_state_field_type_24_is_repeated =
    control_io_metadata_init_bits_desc_state_field_type_24_is_repeated; // @[FpgaCloudSerHw.scala 114:49]
  assign meta_table_io_class_meta_init_bits_desc_state_field_type_24_field_type =
    control_io_metadata_init_bits_desc_state_field_type_24_field_type; // @[FpgaCloudSerHw.scala 114:49]
  assign meta_table_io_class_meta_init_bits_desc_state_field_type_24_sub_class_id =
    control_io_metadata_init_bits_desc_state_field_type_24_sub_class_id; // @[FpgaCloudSerHw.scala 114:49]
  assign meta_table_io_class_meta_init_bits_desc_state_field_type_24_is_host =
    control_io_metadata_init_bits_desc_state_field_type_24_is_host; // @[FpgaCloudSerHw.scala 114:49]
  assign meta_table_io_class_meta_init_bits_desc_state_field_type_25_is_repeated =
    control_io_metadata_init_bits_desc_state_field_type_25_is_repeated; // @[FpgaCloudSerHw.scala 114:49]
  assign meta_table_io_class_meta_init_bits_desc_state_field_type_25_field_type =
    control_io_metadata_init_bits_desc_state_field_type_25_field_type; // @[FpgaCloudSerHw.scala 114:49]
  assign meta_table_io_class_meta_init_bits_desc_state_field_type_25_sub_class_id =
    control_io_metadata_init_bits_desc_state_field_type_25_sub_class_id; // @[FpgaCloudSerHw.scala 114:49]
  assign meta_table_io_class_meta_init_bits_desc_state_field_type_25_is_host =
    control_io_metadata_init_bits_desc_state_field_type_25_is_host; // @[FpgaCloudSerHw.scala 114:49]
  assign meta_table_io_class_meta_init_bits_desc_state_field_type_26_is_repeated =
    control_io_metadata_init_bits_desc_state_field_type_26_is_repeated; // @[FpgaCloudSerHw.scala 114:49]
  assign meta_table_io_class_meta_init_bits_desc_state_field_type_26_field_type =
    control_io_metadata_init_bits_desc_state_field_type_26_field_type; // @[FpgaCloudSerHw.scala 114:49]
  assign meta_table_io_class_meta_init_bits_desc_state_field_type_26_sub_class_id =
    control_io_metadata_init_bits_desc_state_field_type_26_sub_class_id; // @[FpgaCloudSerHw.scala 114:49]
  assign meta_table_io_class_meta_init_bits_desc_state_field_type_26_is_host =
    control_io_metadata_init_bits_desc_state_field_type_26_is_host; // @[FpgaCloudSerHw.scala 114:49]
  assign meta_table_io_class_meta_init_bits_desc_state_field_type_27_is_repeated =
    control_io_metadata_init_bits_desc_state_field_type_27_is_repeated; // @[FpgaCloudSerHw.scala 114:49]
  assign meta_table_io_class_meta_init_bits_desc_state_field_type_27_field_type =
    control_io_metadata_init_bits_desc_state_field_type_27_field_type; // @[FpgaCloudSerHw.scala 114:49]
  assign meta_table_io_class_meta_init_bits_desc_state_field_type_27_sub_class_id =
    control_io_metadata_init_bits_desc_state_field_type_27_sub_class_id; // @[FpgaCloudSerHw.scala 114:49]
  assign meta_table_io_class_meta_init_bits_desc_state_field_type_27_is_host =
    control_io_metadata_init_bits_desc_state_field_type_27_is_host; // @[FpgaCloudSerHw.scala 114:49]
  assign meta_table_io_class_meta_init_bits_desc_state_field_type_28_is_repeated =
    control_io_metadata_init_bits_desc_state_field_type_28_is_repeated; // @[FpgaCloudSerHw.scala 114:49]
  assign meta_table_io_class_meta_init_bits_desc_state_field_type_28_field_type =
    control_io_metadata_init_bits_desc_state_field_type_28_field_type; // @[FpgaCloudSerHw.scala 114:49]
  assign meta_table_io_class_meta_init_bits_desc_state_field_type_28_sub_class_id =
    control_io_metadata_init_bits_desc_state_field_type_28_sub_class_id; // @[FpgaCloudSerHw.scala 114:49]
  assign meta_table_io_class_meta_init_bits_desc_state_field_type_28_is_host =
    control_io_metadata_init_bits_desc_state_field_type_28_is_host; // @[FpgaCloudSerHw.scala 114:49]
  assign meta_table_io_class_meta_init_bits_desc_state_field_type_29_is_repeated =
    control_io_metadata_init_bits_desc_state_field_type_29_is_repeated; // @[FpgaCloudSerHw.scala 114:49]
  assign meta_table_io_class_meta_init_bits_desc_state_field_type_29_field_type =
    control_io_metadata_init_bits_desc_state_field_type_29_field_type; // @[FpgaCloudSerHw.scala 114:49]
  assign meta_table_io_class_meta_init_bits_desc_state_field_type_29_sub_class_id =
    control_io_metadata_init_bits_desc_state_field_type_29_sub_class_id; // @[FpgaCloudSerHw.scala 114:49]
  assign meta_table_io_class_meta_init_bits_desc_state_field_type_29_is_host =
    control_io_metadata_init_bits_desc_state_field_type_29_is_host; // @[FpgaCloudSerHw.scala 114:49]
  assign meta_table_io_class_meta_init_bits_desc_state_field_type_30_is_repeated =
    control_io_metadata_init_bits_desc_state_field_type_30_is_repeated; // @[FpgaCloudSerHw.scala 114:49]
  assign meta_table_io_class_meta_init_bits_desc_state_field_type_30_field_type =
    control_io_metadata_init_bits_desc_state_field_type_30_field_type; // @[FpgaCloudSerHw.scala 114:49]
  assign meta_table_io_class_meta_init_bits_desc_state_field_type_30_sub_class_id =
    control_io_metadata_init_bits_desc_state_field_type_30_sub_class_id; // @[FpgaCloudSerHw.scala 114:49]
  assign meta_table_io_class_meta_init_bits_desc_state_field_type_30_is_host =
    control_io_metadata_init_bits_desc_state_field_type_30_is_host; // @[FpgaCloudSerHw.scala 114:49]
  assign meta_table_io_class_meta_init_bits_desc_state_field_type_31_is_repeated =
    control_io_metadata_init_bits_desc_state_field_type_31_is_repeated; // @[FpgaCloudSerHw.scala 114:49]
  assign meta_table_io_class_meta_init_bits_desc_state_field_type_31_field_type =
    control_io_metadata_init_bits_desc_state_field_type_31_field_type; // @[FpgaCloudSerHw.scala 114:49]
  assign meta_table_io_class_meta_init_bits_desc_state_field_type_31_sub_class_id =
    control_io_metadata_init_bits_desc_state_field_type_31_sub_class_id; // @[FpgaCloudSerHw.scala 114:49]
  assign meta_table_io_class_meta_init_bits_desc_state_field_type_31_is_host =
    control_io_metadata_init_bits_desc_state_field_type_31_is_host; // @[FpgaCloudSerHw.scala 114:49]
  assign meta_table_io_class_meta_init_bits_desc_state_field_type_32_is_repeated =
    control_io_metadata_init_bits_desc_state_field_type_32_is_repeated; // @[FpgaCloudSerHw.scala 114:49]
  assign meta_table_io_class_meta_init_bits_desc_state_field_type_32_field_type =
    control_io_metadata_init_bits_desc_state_field_type_32_field_type; // @[FpgaCloudSerHw.scala 114:49]
  assign meta_table_io_class_meta_init_bits_desc_state_field_type_32_sub_class_id =
    control_io_metadata_init_bits_desc_state_field_type_32_sub_class_id; // @[FpgaCloudSerHw.scala 114:49]
  assign meta_table_io_class_meta_init_bits_desc_state_field_type_32_is_host =
    control_io_metadata_init_bits_desc_state_field_type_32_is_host; // @[FpgaCloudSerHw.scala 114:49]
  assign meta_table_io_s_class_meta_req_valid = ser_io_class_meta_req_valid; // @[FpgaCloudSerHw.scala 121:31]
  assign meta_table_io_s_class_meta_req_bits_class_id = ser_io_class_meta_req_bits_class_id; // @[FpgaCloudSerHw.scala 121:31]
  assign control_clock = clock;
  assign control_reset = ~userRstn; // @[FpgaCloudSerHw.scala 101:33]
  assign control_io_axi_aw_valid = qdma_io_axib_aw_valid; // @[FpgaCloudSerHw.scala 112:57]
  assign control_io_axi_aw_bits_addr = qdma_io_axib_aw_bits_addr; // @[FpgaCloudSerHw.scala 112:57]
  assign control_io_axi_w_valid = qdma_io_axib_w_valid; // @[FpgaCloudSerHw.scala 112:57]
  assign control_io_axi_w_bits_data = qdma_io_axib_w_bits_data; // @[FpgaCloudSerHw.scala 112:57]
  assign control_io_axi_r_ready = qdma_io_axib_r_ready; // @[FpgaCloudSerHw.scala 112:57]
  assign control_io_ser_cmd_ready = ser_io_meta_in_ready; // @[FpgaCloudSerHw.scala 115:49]
  assign instIlaDbg_clk = clock; // @[ILA_VIO.scala 34:25]
  assign instIlaDbg_data_1 = timer_en; // @[ILA_VIO.scala 35:58]
  assign instIlaDbg_data_0 = timer_cnt; // @[ILA_VIO.scala 35:58]
  always @(posedge hbmDriver_io_hbm_clk) begin
    hbmRstn <= hbmDriver_io_hbm_rstn; // @[FpgaCloudSerHw.scala 52:100]
  end
  always @(posedge clock) begin
    if (_T) begin // @[FpgaCloudSerHw.scala 145:39]
      timer_en <= 1'h0; // @[FpgaCloudSerHw.scala 145:39]
    end else begin
      timer_en <= _GEN_1;
    end
    if (_T) begin // @[FpgaCloudSerHw.scala 146:38]
      done_en <= 1'h0; // @[FpgaCloudSerHw.scala 146:38]
    end else if (_T_1) begin // @[FpgaCloudSerHw.scala 172:50]
      done_en <= 1'h0; // @[FpgaCloudSerHw.scala 173:41]
    end else begin
      done_en <= _GEN_4;
    end
    if (_T) begin // @[FpgaCloudSerHw.scala 147:40]
      timer_cnt <= 32'h0; // @[FpgaCloudSerHw.scala 147:40]
    end else if (_T_1) begin // @[FpgaCloudSerHw.scala 157:50]
      timer_cnt <= 32'h0; // @[FpgaCloudSerHw.scala 158:41]
    end else if (timer_en) begin // @[FpgaCloudSerHw.scala 159:38]
      timer_cnt <= _timer_cnt_T_1; // @[FpgaCloudSerHw.scala 160:41]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  hbmRstn = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  timer_en = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  done_en = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  timer_cnt = _RAND_3[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ila_debug(
input clk,
input [31:0] data_0,
input [0:0] data_1);

wire [31:0] timer_cnt = data_0;
wire [0:0] timer_en = data_1;

ila_debug_inner inst_ila_debug(
.clk(clk),
.probe0(timer_cnt), //[31:0]
.probe1(timer_en)); //[0:0]
endmodule
/*
create_ip -name ila -vendor xilinx.com -library ip -version 6.2 -module_name ila_debug_inner
set_property -dict [list CONFIG.C_INPUT_PIPE_STAGES {6} CONFIG.C_PROBE0_WIDTH {32} CONFIG.C_PROBE1_WIDTH {1} CONFIG.C_DATA_DEPTH {1024} CONFIG.C_NUM_OF_PROBES {2} ] [get_ips ila_debug_inner]
*/
