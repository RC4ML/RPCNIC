


`timescale 1ns / 1ns
module tb_cloudfpgaSerSim(

    );

reg                 clock                         =0;
reg                 reset                         =0;
wire                io_axib_aw_ready              ;
reg                 io_axib_aw_valid              =0;
reg       [63:0]    io_axib_aw_bits_addr          =0;
reg       [1:0]     io_axib_aw_bits_burst         =0;
reg       [3:0]     io_axib_aw_bits_cache         =0;
reg       [3:0]     io_axib_aw_bits_id            =0;
reg       [7:0]     io_axib_aw_bits_len           =0;
reg                 io_axib_aw_bits_lock          =0;
reg       [2:0]     io_axib_aw_bits_prot          =0;
reg       [3:0]     io_axib_aw_bits_qos           =0;
reg       [3:0]     io_axib_aw_bits_region        =0;
reg       [2:0]     io_axib_aw_bits_size          =0;
wire                io_axib_ar_ready              ;
reg                 io_axib_ar_valid              =0;
reg       [63:0]    io_axib_ar_bits_addr          =0;
reg       [1:0]     io_axib_ar_bits_burst         =0;
reg       [3:0]     io_axib_ar_bits_cache         =0;
reg       [3:0]     io_axib_ar_bits_id            =0;
reg       [7:0]     io_axib_ar_bits_len           =0;
reg                 io_axib_ar_bits_lock          =0;
reg       [2:0]     io_axib_ar_bits_prot          =0;
reg       [3:0]     io_axib_ar_bits_qos           =0;
reg       [3:0]     io_axib_ar_bits_region        =0;
reg       [2:0]     io_axib_ar_bits_size          =0;
wire                io_axib_w_ready               ;
reg                 io_axib_w_valid               =0;
reg       [511:0]   io_axib_w_bits_data           =0;
reg                 io_axib_w_bits_last           =0;
reg       [63:0]    io_axib_w_bits_strb           =0;
reg                 io_axib_r_ready               =0;
wire                io_axib_r_valid               ;
wire      [511:0]   io_axib_r_bits_data           ;
wire                io_axib_r_bits_last           ;
wire      [1:0]     io_axib_r_bits_resp           ;
wire      [3:0]     io_axib_r_bits_id             ;
reg                 io_axib_b_ready               =0;
wire                io_axib_b_valid               ;
wire      [3:0]     io_axib_b_bits_id             ;
wire      [1:0]     io_axib_b_bits_resp           ;
wire                io_m_mem_read_cmd_ready       ;
wire                io_m_mem_read_cmd_valid       ;
wire      [63:0]    io_m_mem_read_cmd_bits_vaddr  ;
wire      [31:0]    io_m_mem_read_cmd_bits_length ;
wire                io_s_mem_read_data_ready      ;
wire                 io_s_mem_read_data_valid      ;
wire                 io_s_mem_read_data_bits_last  ;
wire       [511:0]   io_s_mem_read_data_bits_data  ;
wire       [63:0]    io_s_mem_read_data_bits_keep  ;
wire                 io_m_mem_write_cmd_ready      ;
wire                io_m_mem_write_cmd_valid      ;
wire      [63:0]    io_m_mem_write_cmd_bits_vaddr ;
wire      [31:0]    io_m_mem_write_cmd_bits_length;
wire                 io_m_mem_write_data_ready     ;
wire                io_m_mem_write_data_valid     ;
wire                io_m_mem_write_data_bits_last ;
wire      [511:0]   io_m_mem_write_data_bits_data ;
wire      [63:0]    io_m_mem_write_data_bits_keep ;
wire      [31:0]    io_status_0                   ;
wire      [31:0]    io_status_1                   ;
wire      [31:0]    io_status_2                   ;
wire      [31:0]    io_status_3                   ;
wire      [31:0]    io_status_4                   ;
wire      [31:0]    io_status_5                   ;
wire      [31:0]    io_status_6                   ;
wire      [31:0]    io_status_7                   ;
wire      [31:0]    io_status_8                   ;
wire      [31:0]    io_status_9                   ;
wire      [31:0]    io_status_10                  ;
wire      [31:0]    io_status_11                  ;
wire      [31:0]    io_status_12                  ;
wire      [31:0]    io_status_13                  ;
wire      [31:0]    io_status_14                  ;
wire      [31:0]    io_status_15                  ;
wire      [31:0]    io_status_16                  ;
wire      [31:0]    io_status_17                  ;
wire      [31:0]    io_status_18                  ;
wire      [31:0]    io_status_19                  ;
wire      [31:0]    io_status_20                  ;
wire      [31:0]    io_status_21                  ;
wire      [31:0]    io_status_22                  ;
wire      [31:0]    io_status_23                  ;
wire      [31:0]    io_status_24                  ;
wire      [31:0]    io_status_25                  ;
wire      [31:0]    io_status_26                  ;
wire      [31:0]    io_status_27                  ;
wire      [31:0]    io_status_28                  ;
wire      [31:0]    io_status_29                  ;
wire      [31:0]    io_status_30                  ;
wire      [31:0]    io_status_31                  ;
wire      [31:0]    io_status_32                  ;
wire      [31:0]    io_status_33                  ;
wire      [31:0]    io_status_34                  ;
wire      [31:0]    io_status_35                  ;
wire      [31:0]    io_status_36                  ;
wire      [31:0]    io_status_37                  ;
wire      [31:0]    io_status_38                  ;
wire      [31:0]    io_status_39                  ;
wire      [31:0]    io_status_40                  ;
wire      [31:0]    io_status_41                  ;
wire      [31:0]    io_status_42                  ;
wire      [31:0]    io_status_43                  ;
wire      [31:0]    io_status_44                  ;
wire      [31:0]    io_status_45                  ;
wire      [31:0]    io_status_46                  ;
wire      [31:0]    io_status_47                  ;
wire      [31:0]    io_status_48                  ;
wire      [31:0]    io_status_49                  ;
wire      [31:0]    io_status_50                  ;
wire      [31:0]    io_status_51                  ;
wire      [31:0]    io_status_52                  ;
wire      [31:0]    io_status_53                  ;
wire      [31:0]    io_status_54                  ;
wire      [31:0]    io_status_55                  ;
wire      [31:0]    io_status_56                  ;
wire      [31:0]    io_status_57                  ;
wire      [31:0]    io_status_58                  ;
wire      [31:0]    io_status_59                  ;
wire      [31:0]    io_status_60                  ;
wire      [31:0]    io_status_61                  ;
wire      [31:0]    io_status_62                  ;
wire      [31:0]    io_status_63                  ;
wire      [31:0]    io_status_64                  ;
wire      [31:0]    io_status_65                  ;
wire      [31:0]    io_status_66                  ;
wire      [31:0]    io_status_67                  ;
wire      [31:0]    io_status_68                  ;
wire      [31:0]    io_status_69                  ;
wire      [31:0]    io_status_70                  ;
wire      [31:0]    io_status_71                  ;
wire      [31:0]    io_status_72                  ;
wire      [31:0]    io_status_73                  ;
wire      [31:0]    io_status_74                  ;
wire      [31:0]    io_status_75                  ;
wire      [31:0]    io_status_76                  ;
wire      [31:0]    io_status_77                  ;
wire      [31:0]    io_status_78                  ;
wire      [31:0]    io_status_79                  ;
wire      [31:0]    io_status_80                  ;
wire      [31:0]    io_status_81                  ;
wire      [31:0]    io_status_82                  ;
wire      [31:0]    io_status_83                  ;
wire      [31:0]    io_status_84                  ;
wire      [31:0]    io_status_85                  ;
wire      [31:0]    io_status_86                  ;
wire      [31:0]    io_status_87                  ;
wire      [31:0]    io_status_88                  ;
wire      [31:0]    io_status_89                  ;
wire      [31:0]    io_status_90                  ;
wire      [31:0]    io_status_91                  ;
wire      [31:0]    io_status_92                  ;
wire      [31:0]    io_status_93                  ;
wire      [31:0]    io_status_94                  ;
wire      [31:0]    io_status_95                  ;
wire      [31:0]    io_status_96                  ;
wire      [31:0]    io_status_97                  ;
wire      [31:0]    io_status_98                  ;
wire      [31:0]    io_status_99                  ;
wire      [31:0]    io_status_100                 ;
wire      [31:0]    io_status_101                 ;
wire      [31:0]    io_status_102                 ;
wire      [31:0]    io_status_103                 ;
wire      [31:0]    io_status_104                 ;
wire      [31:0]    io_status_105                 ;
wire      [31:0]    io_status_106                 ;
wire      [31:0]    io_status_107                 ;
wire      [31:0]    io_status_108                 ;
wire      [31:0]    io_status_109                 ;
wire      [31:0]    io_status_110                 ;
wire      [31:0]    io_status_111                 ;
wire      [31:0]    io_status_112                 ;
wire      [31:0]    io_status_113                 ;
wire      [31:0]    io_status_114                 ;
wire      [31:0]    io_status_115                 ;
wire      [31:0]    io_status_116                 ;
wire      [31:0]    io_status_117                 ;
wire      [31:0]    io_status_118                 ;
wire      [31:0]    io_status_119                 ;
wire      [31:0]    io_status_120                 ;
wire      [31:0]    io_status_121                 ;
wire      [31:0]    io_status_122                 ;
wire      [31:0]    io_status_123                 ;
wire      [31:0]    io_status_124                 ;
wire      [31:0]    io_status_125                 ;
wire      [31:0]    io_status_126                 ;
wire      [31:0]    io_status_127                 ;
wire      [31:0]    io_status_128                 ;
wire      [31:0]    io_status_129                 ;
wire      [31:0]    io_status_130                 ;
wire      [31:0]    io_status_131                 ;
wire      [31:0]    io_status_132                 ;
wire      [31:0]    io_status_133                 ;
wire      [31:0]    io_status_134                 ;
wire      [31:0]    io_status_135                 ;
wire      [31:0]    io_status_136                 ;
wire      [31:0]    io_status_137                 ;
wire      [31:0]    io_status_138                 ;
wire      [31:0]    io_status_139                 ;
wire      [31:0]    io_status_140                 ;
wire      [31:0]    io_status_141                 ;
wire      [31:0]    io_status_142                 ;
wire      [31:0]    io_status_143                 ;
wire      [31:0]    io_status_144                 ;
wire      [31:0]    io_status_145                 ;
wire      [31:0]    io_status_146                 ;
wire      [31:0]    io_status_147                 ;
wire      [31:0]    io_status_148                 ;
wire      [31:0]    io_status_149                 ;
wire      [31:0]    io_status_150                 ;
wire      [31:0]    io_status_151                 ;
wire      [31:0]    io_status_152                 ;
wire      [31:0]    io_status_153                 ;
wire      [31:0]    io_status_154                 ;
wire      [31:0]    io_status_155                 ;
wire      [31:0]    io_status_156                 ;
wire      [31:0]    io_status_157                 ;
wire      [31:0]    io_status_158                 ;
wire      [31:0]    io_status_159                 ;
wire      [31:0]    io_status_160                 ;
wire      [31:0]    io_status_161                 ;
wire      [31:0]    io_status_162                 ;
wire      [31:0]    io_status_163                 ;
wire      [31:0]    io_status_164                 ;
wire      [31:0]    io_status_165                 ;
wire      [31:0]    io_status_166                 ;
wire      [31:0]    io_status_167                 ;
wire      [31:0]    io_status_168                 ;
wire      [31:0]    io_status_169                 ;
wire      [31:0]    io_status_170                 ;
wire      [31:0]    io_status_171                 ;
wire      [31:0]    io_status_172                 ;
wire      [31:0]    io_status_173                 ;
wire      [31:0]    io_status_174                 ;
wire      [31:0]    io_status_175                 ;
wire      [31:0]    io_status_176                 ;
wire      [31:0]    io_status_177                 ;
wire      [31:0]    io_status_178                 ;
wire      [31:0]    io_status_179                 ;
wire      [31:0]    io_status_180                 ;
wire      [31:0]    io_status_181                 ;
wire      [31:0]    io_status_182                 ;
wire      [31:0]    io_status_183                 ;
wire      [31:0]    io_status_184                 ;
wire      [31:0]    io_status_185                 ;
wire      [31:0]    io_status_186                 ;
wire      [31:0]    io_status_187                 ;
wire      [31:0]    io_status_188                 ;
wire      [31:0]    io_status_189                 ;
wire      [31:0]    io_status_190                 ;
wire      [31:0]    io_status_191                 ;
wire      [31:0]    io_status_192                 ;
wire      [31:0]    io_status_193                 ;
wire      [31:0]    io_status_194                 ;
wire      [31:0]    io_status_195                 ;
wire      [31:0]    io_status_196                 ;
wire      [31:0]    io_status_197                 ;
wire      [31:0]    io_status_198                 ;
wire      [31:0]    io_status_199                 ;
wire      [31:0]    io_status_200                 ;
wire      [31:0]    io_status_201                 ;
wire      [31:0]    io_status_202                 ;
wire      [31:0]    io_status_203                 ;
wire      [31:0]    io_status_204                 ;
wire      [31:0]    io_status_205                 ;
wire      [31:0]    io_status_206                 ;
wire      [31:0]    io_status_207                 ;
wire      [31:0]    io_status_208                 ;
wire      [31:0]    io_status_209                 ;
wire      [31:0]    io_status_210                 ;
wire      [31:0]    io_status_211                 ;
wire      [31:0]    io_status_212                 ;
wire      [31:0]    io_status_213                 ;
wire      [31:0]    io_status_214                 ;
wire      [31:0]    io_status_215                 ;
wire      [31:0]    io_status_216                 ;
wire      [31:0]    io_status_217                 ;
wire      [31:0]    io_status_218                 ;
wire      [31:0]    io_status_219                 ;
wire      [31:0]    io_status_220                 ;
wire      [31:0]    io_status_221                 ;
wire      [31:0]    io_status_222                 ;
wire      [31:0]    io_status_223                 ;
wire      [31:0]    io_status_224                 ;
wire      [31:0]    io_status_225                 ;
wire      [31:0]    io_status_226                 ;
wire      [31:0]    io_status_227                 ;
wire      [31:0]    io_status_228                 ;
wire      [31:0]    io_status_229                 ;
wire      [31:0]    io_status_230                 ;
wire      [31:0]    io_status_231                 ;
wire      [31:0]    io_status_232                 ;
wire      [31:0]    io_status_233                 ;
wire      [31:0]    io_status_234                 ;
wire      [31:0]    io_status_235                 ;
wire      [31:0]    io_status_236                 ;
wire      [31:0]    io_status_237                 ;
wire      [31:0]    io_status_238                 ;
wire      [31:0]    io_status_239                 ;
wire      [31:0]    io_status_240                 ;
wire      [31:0]    io_status_241                 ;
wire      [31:0]    io_status_242                 ;
wire      [31:0]    io_status_243                 ;
wire      [31:0]    io_status_244                 ;
wire      [31:0]    io_status_245                 ;
wire      [31:0]    io_status_246                 ;
wire      [31:0]    io_status_247                 ;
wire      [31:0]    io_status_248                 ;
wire      [31:0]    io_status_249                 ;
wire      [31:0]    io_status_250                 ;
wire      [31:0]    io_status_251                 ;
wire      [31:0]    io_status_252                 ;
wire      [31:0]    io_status_253                 ;
wire      [31:0]    io_status_254                 ;
wire      [31:0]    io_status_255                 ;
wire      [31:0]    io_status_256                 ;
wire      [31:0]    io_status_257                 ;
wire      [31:0]    io_status_258                 ;
wire      [31:0]    io_status_259                 ;
wire      [31:0]    io_status_260                 ;
wire      [31:0]    io_status_261                 ;
wire      [31:0]    io_status_262                 ;
wire      [31:0]    io_status_263                 ;
wire      [31:0]    io_status_264                 ;
wire      [31:0]    io_status_265                 ;
wire      [31:0]    io_status_266                 ;
wire      [31:0]    io_status_267                 ;
wire      [31:0]    io_status_268                 ;
wire      [31:0]    io_status_269                 ;
wire      [31:0]    io_status_270                 ;
wire      [31:0]    io_status_271                 ;
wire      [31:0]    io_status_272                 ;
wire      [31:0]    io_status_273                 ;
wire      [31:0]    io_status_274                 ;
wire      [31:0]    io_status_275                 ;
wire      [31:0]    io_status_276                 ;
wire      [31:0]    io_status_277                 ;
wire      [31:0]    io_status_278                 ;
wire      [31:0]    io_status_279                 ;
wire      [31:0]    io_status_280                 ;
wire      [31:0]    io_status_281                 ;
wire      [31:0]    io_status_282                 ;
wire      [31:0]    io_status_283                 ;
wire      [31:0]    io_status_284                 ;
wire      [31:0]    io_status_285                 ;
wire      [31:0]    io_status_286                 ;
wire      [31:0]    io_status_287                 ;
wire      [31:0]    io_status_288                 ;
wire      [31:0]    io_status_289                 ;
wire      [31:0]    io_status_290                 ;
wire      [31:0]    io_status_291                 ;
wire      [31:0]    io_status_292                 ;
wire      [31:0]    io_status_293                 ;
wire      [31:0]    io_status_294                 ;
wire      [31:0]    io_status_295                 ;
wire      [31:0]    io_status_296                 ;
wire      [31:0]    io_status_297                 ;
wire      [31:0]    io_status_298                 ;
wire      [31:0]    io_status_299                 ;
wire      [31:0]    io_status_300                 ;
wire      [31:0]    io_status_301                 ;
wire      [31:0]    io_status_302                 ;
wire      [31:0]    io_status_303                 ;
wire      [31:0]    io_status_304                 ;
wire      [31:0]    io_status_305                 ;
wire      [31:0]    io_status_306                 ;
wire      [31:0]    io_status_307                 ;
wire      [31:0]    io_status_308                 ;
wire      [31:0]    io_status_309                 ;
wire      [31:0]    io_status_310                 ;
wire      [31:0]    io_status_311                 ;
wire      [31:0]    io_status_312                 ;
wire      [31:0]    io_status_313                 ;
wire      [31:0]    io_status_314                 ;
wire      [31:0]    io_status_315                 ;
wire      [31:0]    io_status_316                 ;
wire      [31:0]    io_status_317                 ;
wire      [31:0]    io_status_318                 ;
wire      [31:0]    io_status_319                 ;
wire      [31:0]    io_status_320                 ;
wire      [31:0]    io_status_321                 ;
wire      [31:0]    io_status_322                 ;
wire      [31:0]    io_status_323                 ;
wire      [31:0]    io_status_324                 ;
wire      [31:0]    io_status_325                 ;
wire      [31:0]    io_status_326                 ;
wire      [31:0]    io_status_327                 ;
wire      [31:0]    io_status_328                 ;
wire      [31:0]    io_status_329                 ;
wire      [31:0]    io_status_330                 ;
wire      [31:0]    io_status_331                 ;
wire      [31:0]    io_status_332                 ;
wire      [31:0]    io_status_333                 ;
wire      [31:0]    io_status_334                 ;
wire      [31:0]    io_status_335                 ;
wire      [31:0]    io_status_336                 ;
wire      [31:0]    io_status_337                 ;
wire      [31:0]    io_status_338                 ;
wire      [31:0]    io_status_339                 ;
wire      [31:0]    io_status_340                 ;
wire      [31:0]    io_status_341                 ;
wire      [31:0]    io_status_342                 ;
wire      [31:0]    io_status_343                 ;
wire      [31:0]    io_status_344                 ;
wire      [31:0]    io_status_345                 ;
wire      [31:0]    io_status_346                 ;
wire      [31:0]    io_status_347                 ;
wire      [31:0]    io_status_348                 ;
wire      [31:0]    io_status_349                 ;
wire      [31:0]    io_status_350                 ;
wire      [31:0]    io_status_351                 ;
wire      [31:0]    io_status_352                 ;
wire      [31:0]    io_status_353                 ;
wire      [31:0]    io_status_354                 ;
wire      [31:0]    io_status_355                 ;
wire      [31:0]    io_status_356                 ;
wire      [31:0]    io_status_357                 ;
wire      [31:0]    io_status_358                 ;
wire      [31:0]    io_status_359                 ;
wire      [31:0]    io_status_360                 ;
wire      [31:0]    io_status_361                 ;
wire      [31:0]    io_status_362                 ;
wire      [31:0]    io_status_363                 ;
wire      [31:0]    io_status_364                 ;
wire      [31:0]    io_status_365                 ;
wire      [31:0]    io_status_366                 ;
wire      [31:0]    io_status_367                 ;
wire      [31:0]    io_status_368                 ;
wire      [31:0]    io_status_369                 ;
wire      [31:0]    io_status_370                 ;
wire      [31:0]    io_status_371                 ;
wire      [31:0]    io_status_372                 ;
wire      [31:0]    io_status_373                 ;
wire      [31:0]    io_status_374                 ;
wire      [31:0]    io_status_375                 ;
wire      [31:0]    io_status_376                 ;
wire      [31:0]    io_status_377                 ;
wire      [31:0]    io_status_378                 ;
wire      [31:0]    io_status_379                 ;
wire      [31:0]    io_status_380                 ;
wire      [31:0]    io_status_381                 ;
wire      [31:0]    io_status_382                 ;
wire      [31:0]    io_status_383                 ;
wire      [31:0]    io_status_384                 ;
wire      [31:0]    io_status_385                 ;
wire      [31:0]    io_status_386                 ;
wire      [31:0]    io_status_387                 ;
wire      [31:0]    io_status_388                 ;
wire      [31:0]    io_status_389                 ;
wire      [31:0]    io_status_390                 ;
wire      [31:0]    io_status_391                 ;
wire      [31:0]    io_status_392                 ;
wire      [31:0]    io_status_393                 ;
wire      [31:0]    io_status_394                 ;
wire      [31:0]    io_status_395                 ;
wire      [31:0]    io_status_396                 ;
wire      [31:0]    io_status_397                 ;
wire      [31:0]    io_status_398                 ;
wire      [31:0]    io_status_399                 ;
wire      [31:0]    io_status_400                 ;
wire      [31:0]    io_status_401                 ;
wire      [31:0]    io_status_402                 ;
wire      [31:0]    io_status_403                 ;
wire      [31:0]    io_status_404                 ;
wire      [31:0]    io_status_405                 ;
wire      [31:0]    io_status_406                 ;
wire      [31:0]    io_status_407                 ;
wire      [31:0]    io_status_408                 ;
wire      [31:0]    io_status_409                 ;
wire      [31:0]    io_status_410                 ;
wire      [31:0]    io_status_411                 ;
wire      [31:0]    io_status_412                 ;
wire      [31:0]    io_status_413                 ;
wire      [31:0]    io_status_414                 ;
wire      [31:0]    io_status_415                 ;
wire      [31:0]    io_status_416                 ;
wire      [31:0]    io_status_417                 ;
wire      [31:0]    io_status_418                 ;
wire      [31:0]    io_status_419                 ;
wire      [31:0]    io_status_420                 ;
wire      [31:0]    io_status_421                 ;
wire      [31:0]    io_status_422                 ;
wire      [31:0]    io_status_423                 ;
wire      [31:0]    io_status_424                 ;
wire      [31:0]    io_status_425                 ;
wire      [31:0]    io_status_426                 ;
wire      [31:0]    io_status_427                 ;
wire      [31:0]    io_status_428                 ;
wire      [31:0]    io_status_429                 ;
wire      [31:0]    io_status_430                 ;
wire      [31:0]    io_status_431                 ;
wire      [31:0]    io_status_432                 ;
wire      [31:0]    io_status_433                 ;
wire      [31:0]    io_status_434                 ;
wire      [31:0]    io_status_435                 ;
wire      [31:0]    io_status_436                 ;
wire      [31:0]    io_status_437                 ;
wire      [31:0]    io_status_438                 ;
wire      [31:0]    io_status_439                 ;
wire      [31:0]    io_status_440                 ;
wire      [31:0]    io_status_441                 ;
wire      [31:0]    io_status_442                 ;
wire      [31:0]    io_status_443                 ;
wire      [31:0]    io_status_444                 ;
wire      [31:0]    io_status_445                 ;
wire      [31:0]    io_status_446                 ;
wire      [31:0]    io_status_447                 ;
wire      [31:0]    io_status_448                 ;
wire      [31:0]    io_status_449                 ;
wire      [31:0]    io_status_450                 ;
wire      [31:0]    io_status_451                 ;
wire      [31:0]    io_status_452                 ;
wire      [31:0]    io_status_453                 ;
wire      [31:0]    io_status_454                 ;
wire      [31:0]    io_status_455                 ;
wire      [31:0]    io_status_456                 ;
wire      [31:0]    io_status_457                 ;
wire      [31:0]    io_status_458                 ;
wire      [31:0]    io_status_459                 ;
wire      [31:0]    io_status_460                 ;
wire      [31:0]    io_status_461                 ;
wire      [31:0]    io_status_462                 ;
wire      [31:0]    io_status_463                 ;
wire      [31:0]    io_status_464                 ;
wire      [31:0]    io_status_465                 ;
wire      [31:0]    io_status_466                 ;
wire      [31:0]    io_status_467                 ;
wire      [31:0]    io_status_468                 ;
wire      [31:0]    io_status_469                 ;
wire      [31:0]    io_status_470                 ;
wire      [31:0]    io_status_471                 ;
wire      [31:0]    io_status_472                 ;
wire      [31:0]    io_status_473                 ;
wire      [31:0]    io_status_474                 ;
wire      [31:0]    io_status_475                 ;
wire      [31:0]    io_status_476                 ;
wire      [31:0]    io_status_477                 ;
wire      [31:0]    io_status_478                 ;
wire      [31:0]    io_status_479                 ;
wire      [31:0]    io_status_480                 ;
wire      [31:0]    io_status_481                 ;
wire      [31:0]    io_status_482                 ;
wire      [31:0]    io_status_483                 ;
wire      [31:0]    io_status_484                 ;
wire      [31:0]    io_status_485                 ;
wire      [31:0]    io_status_486                 ;
wire      [31:0]    io_status_487                 ;
wire      [31:0]    io_status_488                 ;
wire      [31:0]    io_status_489                 ;
wire      [31:0]    io_status_490                 ;
wire      [31:0]    io_status_491                 ;
wire      [31:0]    io_status_492                 ;
wire      [31:0]    io_status_493                 ;
wire      [31:0]    io_status_494                 ;
wire      [31:0]    io_status_495                 ;
wire      [31:0]    io_status_496                 ;
wire      [31:0]    io_status_497                 ;
wire      [31:0]    io_status_498                 ;
wire      [31:0]    io_status_499                 ;
wire      [31:0]    io_status_500                 ;
wire      [31:0]    io_status_501                 ;
wire      [31:0]    io_status_502                 ;
wire      [31:0]    io_status_503                 ;
wire      [31:0]    io_status_504                 ;
wire      [31:0]    io_status_505                 ;
wire      [31:0]    io_status_506                 ;
wire      [31:0]    io_status_507                 ;
wire      [31:0]    io_status_508                 ;
wire      [31:0]    io_status_509                 ;
wire      [31:0]    io_status_510                 ;
wire      [31:0]    io_status_511                 ;



IN#(97)in_io_axib_aw(
        clock,
        reset,
        {io_axib_aw_bits_addr,io_axib_aw_bits_burst,io_axib_aw_bits_cache,io_axib_aw_bits_id,io_axib_aw_bits_len,io_axib_aw_bits_lock,io_axib_aw_bits_prot,io_axib_aw_bits_qos,io_axib_aw_bits_region,io_axib_aw_bits_size},
        io_axib_aw_valid,
        io_axib_aw_ready
);
// addr, burst, cache, id, len, lock, prot, qos, region, size
// 64'h0, 2'h0, 4'h0, 4'h0, 8'h0, 1'h0, 3'h0, 4'h0, 4'h0, 3'h0

IN#(97)in_io_axib_ar(
        clock,
        reset,
        {io_axib_ar_bits_addr,io_axib_ar_bits_burst,io_axib_ar_bits_cache,io_axib_ar_bits_id,io_axib_ar_bits_len,io_axib_ar_bits_lock,io_axib_ar_bits_prot,io_axib_ar_bits_qos,io_axib_ar_bits_region,io_axib_ar_bits_size},
        io_axib_ar_valid,
        io_axib_ar_ready
);
// addr, burst, cache, id, len, lock, prot, qos, region, size
// 64'h0, 2'h0, 4'h0, 4'h0, 8'h0, 1'h0, 3'h0, 4'h0, 4'h0, 3'h0

IN#(577)in_io_axib_w(
        clock,
        reset,
        {io_axib_w_bits_data,io_axib_w_bits_last,io_axib_w_bits_strb},
        io_axib_w_valid,
        io_axib_w_ready
);
// data, last, strb
// 512'h0, 1'h0, 64'h0

OUT#(519)out_io_axib_r(
        clock,
        reset,
        {io_axib_r_bits_data,io_axib_r_bits_last,io_axib_r_bits_resp,io_axib_r_bits_id},
        io_axib_r_valid,
        io_axib_r_ready
);
// data, last, resp, id
// 512'h0, 1'h0, 2'h0, 4'h0

OUT#(6)out_io_axib_b(
        clock,
        reset,
        {io_axib_b_bits_id,io_axib_b_bits_resp},
        io_axib_b_valid,
        io_axib_b_ready
);
// id, resp
// 4'h0, 2'h0





DMA #(512) qdma(
    clock,
    reset,
    //DMA CMD streams
    io_m_mem_read_cmd_valid,
    io_m_mem_read_cmd_ready,
    io_m_mem_read_cmd_bits_vaddr,
    io_m_mem_read_cmd_bits_length,
    io_m_mem_write_cmd_valid,
    io_m_mem_write_cmd_ready,
    io_m_mem_write_cmd_bits_vaddr,
    io_m_mem_write_cmd_bits_length,        
    //DMA Data streams      
    io_s_mem_read_data_valid,
    io_s_mem_read_data_ready,
    io_s_mem_read_data_bits_data,
    io_s_mem_read_data_bits_keep,
    io_s_mem_read_data_bits_last,
    io_m_mem_write_data_valid,
    io_m_mem_write_data_ready,
    io_m_mem_write_data_bits_data,
    io_m_mem_write_data_bits_keep,
    io_m_mem_write_data_bits_last        
);





cloudfpgaSerSim cloudfpgaSerSim_inst(
        .*
);

/*
addr,burst,cache,id,len,lock,prot,qos,region,size
in_io_axib_aw.write({64'h0,2'h0,4'h0,4'h0,8'h0,1'h0,3'h0,4'h0,4'h0,3'h0});

addr,burst,cache,id,len,lock,prot,qos,region,size
in_io_axib_ar.write({64'h0,2'h0,4'h0,4'h0,8'h0,1'h0,3'h0,4'h0,4'h0,3'h0});

data,last,strb
in_io_axib_w.write({512'h0,1'h0,64'h0});

last,data,keep
in_io_s_mem_read_data.write({1'h0,512'h0,64'h0});

*/

reg [511:0] meta_fifo[90:0];
// reg [511:0] h_fifo[1:0];
integer i,j;

initial begin
        reset <= 1;
        clock = 1;
        // $readmemh("/home/amax/hhj/cloud_fpga/serialization/tb/device.txt",d_fifo,0,5);
        $readmemh("/home/amax/hhj/cloud_fpga/cloud_fpga/tb/meta0.txt",meta_fifo,0,90);        
        #1000;
        reset <= 0;
        #100;
        out_io_axib_r.start();
        out_io_axib_b.start();

        for(i=0;i<30;i++) begin
                in_io_axib_aw.write({64'h500,2'h0,4'h0,4'h0,8'h0,1'h0,3'h0,4'h0,4'h0,3'h0});
                in_io_axib_w.write({meta_fifo[i*3],1'h0,64'h0});
                in_io_axib_aw.write({64'h540,2'h0,4'h0,4'h0,8'h0,1'h0,3'h0,4'h0,4'h0,3'h0});
                in_io_axib_w.write({meta_fifo[i*3+1],1'h0,64'h0});
                in_io_axib_aw.write({64'h580,2'h0,4'h0,4'h0,8'h0,1'h0,3'h0,4'h0,4'h0,3'h0});
                in_io_axib_w.write({meta_fifo[i*3+2],1'h0,64'h0});
                #100;
        end


        // in_io_metadata_init.write({10'd1,16'd0,8'd9,1'd0,5'd0,10'd0,1'd0,1'd0,5'd5,10'd0,1'd1,1'd0,5'd3,10'd0,1'd1,1'd0,5'd1,10'd0,1'd0,1'd0,5'd2,10'd0,1'd0,1'd0,5'd6,10'd0,1'd0,1'd0,5'd7,10'd0,1'd1,1'd0,5'd9,10'd0,1'd1,1'd0,5'd11,10'd2,1'd1,1'd1,5'd5,10'd0,1'd1,1'd0,5'd0,10'd0,1'd0,1'd0,5'd0,10'd0,1'd0,1'd0,5'd0,10'd0,1'd0,1'd0,5'd0,10'd0,1'd0,1'd0,5'd0,10'd0,1'd0,1'd0,5'd0,10'd0,1'd0,1'h0,5'h0,10'h0,1'h0,1'h0,5'h0,10'h0,1'h0,1'h0,5'h0,10'h0,1'h0,1'h0,5'h0,10'h0,1'h0,1'h0,5'h0,10'h0,1'h0,1'h0,5'h0,10'h0,1'h0,1'h0,5'h0,10'h0,1'h0,1'h0,5'h0,10'h0,1'h0,1'h0,5'h0,10'h0,1'h0,1'h0,5'h0,10'h0,1'h0,1'h0,5'h0,10'h0,1'h0,1'h0,5'h0,10'h0,1'h0,1'h0,5'h0,10'h0,1'h0,1'h0,5'h0,10'h0,1'h0,1'h0,5'h0,10'h0,1'h0,1'h0,5'h0,10'h0,1'h0,1'h0,5'h0,10'h0,1'h0,1'h0,5'h0,10'h0,1'h0,1'h0,5'h0,10'h0,1'h0,1'h0,5'h0,10'h0,1'h0,1'h0,5'h0,10'h0,1'h0,1'h0,5'h0,10'h0,1'h0,1'h0,5'h0,10'h0,1'h0,1'h0,5'h0,10'h0,1'h0,1'h0,5'h0,10'h0,1'h0,1'h0,5'h0,10'h0,1'h0,1'h0,5'h0,10'h0,1'h0,1'h0,5'h0,10'h0,1'h0,1'h0,5'h0,10'h0,1'h0,1'h0,5'h0,10'h0,1'h0,1'h0,5'h0,10'h0,1'h0,1'h0,5'h0,10'h0,1'h0});
        // in_io_metadata_init.write({10'd2,16'd0,8'd2,1'd0,5'd0,10'd0,1'd0,1'd0,5'd5,10'd0,1'd1,1'd0,5'd9,10'd0,1'd0,1'd0,5'd0,10'd0,1'd0,1'd0,5'd0,10'd0,1'd0,1'd0,5'd0,10'd0,1'd0,1'd0,5'd0,10'd0,1'd0,1'd0,5'd0,10'd0,1'd0,1'd0,5'd0,10'd0,1'd0,1'd0,5'd0,10'd0,1'd0,1'd0,5'd0,10'd0,1'd0,1'd0,5'd0,10'd0,1'd0,1'd0,5'd0,10'd0,1'd0,1'd0,5'd0,10'd0,1'd0,1'd0,5'd0,10'd0,1'd0,1'd0,5'd0,10'd0,1'd0,1'h0,5'h0,10'h0,1'h0,1'h0,5'h0,10'h0,1'h0,1'h0,5'h0,10'h0,1'h0,1'h0,5'h0,10'h0,1'h0,1'h0,5'h0,10'h0,1'h0,1'h0,5'h0,10'h0,1'h0,1'h0,5'h0,10'h0,1'h0,1'h0,5'h0,10'h0,1'h0,1'h0,5'h0,10'h0,1'h0,1'h0,5'h0,10'h0,1'h0,1'h0,5'h0,10'h0,1'h0,1'h0,5'h0,10'h0,1'h0,1'h0,5'h0,10'h0,1'h0,1'h0,5'h0,10'h0,1'h0,1'h0,5'h0,10'h0,1'h0,1'h0,5'h0,10'h0,1'h0,1'h0,5'h0,10'h0,1'h0,1'h0,5'h0,10'h0,1'h0,1'h0,5'h0,10'h0,1'h0,1'h0,5'h0,10'h0,1'h0,1'h0,5'h0,10'h0,1'h0,1'h0,5'h0,10'h0,1'h0,1'h0,5'h0,10'h0,1'h0,1'h0,5'h0,10'h0,1'h0,1'h0,5'h0,10'h0,1'h0,1'h0,5'h0,10'h0,1'h0,1'h0,5'h0,10'h0,1'h0,1'h0,5'h0,10'h0,1'h0,1'h0,5'h0,10'h0,1'h0,1'h0,5'h0,10'h0,1'h0,1'h0,5'h0,10'h0,1'h0,1'h0,5'h0,10'h0,1'h0});    
        qdma.init_from_file("/home/amax/hhj/cloud_fpga/cloud_fpga/tb/rpc0.txt");
        #50;
        in_io_axib_aw.write({64'h340,2'h0,4'h0,4'h0,8'h0,1'h0,3'h0,4'h0,4'h0,3'h0});
        in_io_axib_w.write({512'h2_00000000_00000000_00000000_00000480_0007ee40_00000000,1'h0,64'h0});
        #20000;
        in_io_axib_aw.write({64'h300,2'h0,4'h0,4'h0,8'h0,1'h0,3'h0,4'h0,4'h0,3'h0});
        in_io_axib_w.write({512'h1000_0007ee40_00000447_00000000_00000000_00000000_00000000_00000000_00000119,1'h0,64'h0});

        // in_io_ser_cmd.write({10'h1,32'd35,32'h180,64'h0,64'h0,16'h100});


end

always #5 clock=~clock;
endmodule